// nios_system.v

// Generated using ACDS version 17.1 593

`timescale 1 ps / 1 ps
module nios_system (
		inout  wire        audio_and_video_config_external_interface_SDAT, // audio_and_video_config_external_interface.SDAT
		output wire        audio_and_video_config_external_interface_SCLK, //                                          .SCLK
		output wire        audio_clk_out_clk,                              //                             audio_clk_out.clk
		input  wire        audio_external_interface_ADCDAT,                //                  audio_external_interface.ADCDAT
		input  wire        audio_external_interface_ADCLRCK,               //                                          .ADCLRCK
		input  wire        audio_external_interface_BCLK,                  //                                          .BCLK
		output wire        audio_external_interface_DACDAT,                //                                          .DACDAT
		input  wire        audio_external_interface_DACLRCK,               //                                          .DACLRCK
		inout  wire [7:0]  char_lcd_external_interface_DATA,               //               char_lcd_external_interface.DATA
		output wire        char_lcd_external_interface_ON,                 //                                          .ON
		output wire        char_lcd_external_interface_BLON,               //                                          .BLON
		output wire        char_lcd_external_interface_EN,                 //                                          .EN
		output wire        char_lcd_external_interface_RS,                 //                                          .RS
		output wire        char_lcd_external_interface_RW,                 //                                          .RW
		input  wire        clk_50_2_in_clk,                                //                               clk_50_2_in.clk
		input  wire        clk_50_3_in_clk,                                //                               clk_50_3_in.clk
		input  wire        clk_50_in_clk,                                  //                                 clk_50_in.clk
		output wire [22:0] flash_bridge_out_tcm_address_out,               //                          flash_bridge_out.tcm_address_out
		output wire [0:0]  flash_bridge_out_tcm_read_n_out,                //                                          .tcm_read_n_out
		output wire [0:0]  flash_bridge_out_tcm_write_n_out,               //                                          .tcm_write_n_out
		inout  wire [7:0]  flash_bridge_out_tcm_data_out,                  //                                          .tcm_data_out
		output wire [0:0]  flash_bridge_out_tcm_chipselect_n_out,          //                                          .tcm_chipselect_n_out
		output wire [8:0]  green_led_external_interface_export,            //              green_led_external_interface.export
		output wire [6:0]  hex3_hex0_external_interface_HEX0,              //              hex3_hex0_external_interface.HEX0
		output wire [6:0]  hex3_hex0_external_interface_HEX1,              //                                          .HEX1
		output wire [6:0]  hex3_hex0_external_interface_HEX2,              //                                          .HEX2
		output wire [6:0]  hex3_hex0_external_interface_HEX3,              //                                          .HEX3
		output wire [6:0]  hex7_hex4_external_interface_HEX4,              //              hex7_hex4_external_interface.HEX4
		output wire [6:0]  hex7_hex4_external_interface_HEX5,              //                                          .HEX5
		output wire [6:0]  hex7_hex4_external_interface_HEX6,              //                                          .HEX6
		output wire [6:0]  hex7_hex4_external_interface_HEX7,              //                                          .HEX7
		output wire        mtl_clk_out_clk,                                //                               mtl_clk_out.clk
		output wire        mtl_controller_external_interface_CLK,          //         mtl_controller_external_interface.CLK
		output wire        mtl_controller_external_interface_HS,           //                                          .HS
		output wire        mtl_controller_external_interface_VS,           //                                          .VS
		output wire        mtl_controller_external_interface_DATA_EN,      //                                          .DATA_EN
		output wire [7:0]  mtl_controller_external_interface_R,            //                                          .R
		output wire [7:0]  mtl_controller_external_interface_G,            //                                          .G
		output wire [7:0]  mtl_controller_external_interface_B,            //                                          .B
		inout  wire        ps2_key_external_interface_CLK,                 //                ps2_key_external_interface.CLK
		inout  wire        ps2_key_external_interface_DAT,                 //                                          .DAT
		inout  wire        ps2_mouse_external_interface_CLK,               //              ps2_mouse_external_interface.CLK
		inout  wire        ps2_mouse_external_interface_DAT,               //                                          .DAT
		input  wire [3:0]  pushbuttons_external_interface_export,          //            pushbuttons_external_interface.export
		output wire [17:0] red_leds_external_interface_export,             //               red_leds_external_interface.export
		input  wire        reset_bridge_in_reset_n,                        //                           reset_bridge_in.reset_n
		inout  wire        sd_card_conduit_end_b_SD_cmd,                   //                       sd_card_conduit_end.b_SD_cmd
		inout  wire        sd_card_conduit_end_b_SD_dat,                   //                                          .b_SD_dat
		inout  wire        sd_card_conduit_end_b_SD_dat3,                  //                                          .b_SD_dat3
		output wire        sd_card_conduit_end_o_SD_clock,                 //                                          .o_SD_clock
		output wire        sdram_clk_out_clk,                              //                             sdram_clk_out.clk
		output wire [12:0] sdram_wire_addr,                                //                                sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                                  //                                          .ba
		output wire        sdram_wire_cas_n,                               //                                          .cas_n
		output wire        sdram_wire_cke,                                 //                                          .cke
		output wire        sdram_wire_cs_n,                                //                                          .cs_n
		inout  wire [31:0] sdram_wire_dq,                                  //                                          .dq
		output wire [3:0]  sdram_wire_dqm,                                 //                                          .dqm
		output wire        sdram_wire_ras_n,                               //                                          .ras_n
		output wire        sdram_wire_we_n,                                //                                          .we_n
		input  wire        serial_port_external_interface_RXD,             //            serial_port_external_interface.RXD
		output wire        serial_port_external_interface_TXD,             //                                          .TXD
		inout  wire [15:0] sram_external_interface_DQ,                     //                   sram_external_interface.DQ
		output wire [19:0] sram_external_interface_ADDR,                   //                                          .ADDR
		output wire        sram_external_interface_LB_N,                   //                                          .LB_N
		output wire        sram_external_interface_UB_N,                   //                                          .UB_N
		output wire        sram_external_interface_CE_N,                   //                                          .CE_N
		output wire        sram_external_interface_OE_N,                   //                                          .OE_N
		output wire        sram_external_interface_WE_N,                   //                                          .WE_N
		input  wire [17:0] switches_external_interface_export,             //               switches_external_interface.export
		output wire        sys_clk_out_clk,                                //                               sys_clk_out.clk
		input  wire        video_decoder_external_interface_TD_CLK27,      //          video_decoder_external_interface.TD_CLK27
		input  wire [7:0]  video_decoder_external_interface_TD_DATA,       //                                          .TD_DATA
		input  wire        video_decoder_external_interface_TD_HS,         //                                          .TD_HS
		input  wire        video_decoder_external_interface_TD_VS,         //                                          .TD_VS
		input  wire        video_decoder_external_interface_clk27_reset,   //                                          .clk27_reset
		output wire        video_decoder_external_interface_TD_RESET,      //                                          .TD_RESET
		output wire        video_decoder_external_interface_overflow_flag  //                                          .overflow_flag
	);

	wire         alpha_blending_avalon_blended_source_valid;                                        // alpha_blending:output_valid -> mtl_dual_clock_buffer:stream_in_valid
	wire  [29:0] alpha_blending_avalon_blended_source_data;                                         // alpha_blending:output_data -> mtl_dual_clock_buffer:stream_in_data
	wire         alpha_blending_avalon_blended_source_ready;                                        // mtl_dual_clock_buffer:stream_in_ready -> alpha_blending:output_ready
	wire         alpha_blending_avalon_blended_source_startofpacket;                                // alpha_blending:output_startofpacket -> mtl_dual_clock_buffer:stream_in_startofpacket
	wire         alpha_blending_avalon_blended_source_endofpacket;                                  // alpha_blending:output_endofpacket -> mtl_dual_clock_buffer:stream_in_endofpacket
	wire         mtl_char_buffer_avalon_char_source_valid;                                          // mtl_char_buffer:stream_valid -> alpha_blending:foreground_valid
	wire  [39:0] mtl_char_buffer_avalon_char_source_data;                                           // mtl_char_buffer:stream_data -> alpha_blending:foreground_data
	wire         mtl_char_buffer_avalon_char_source_ready;                                          // alpha_blending:foreground_ready -> mtl_char_buffer:stream_ready
	wire         mtl_char_buffer_avalon_char_source_startofpacket;                                  // mtl_char_buffer:stream_startofpacket -> alpha_blending:foreground_startofpacket
	wire         mtl_char_buffer_avalon_char_source_endofpacket;                                    // mtl_char_buffer:stream_endofpacket -> alpha_blending:foreground_endofpacket
	wire         video_chroma_resampler_avalon_chroma_source_valid;                                 // video_chroma_resampler:stream_out_valid -> video_csc:stream_in_valid
	wire  [23:0] video_chroma_resampler_avalon_chroma_source_data;                                  // video_chroma_resampler:stream_out_data -> video_csc:stream_in_data
	wire         video_chroma_resampler_avalon_chroma_source_ready;                                 // video_csc:stream_in_ready -> video_chroma_resampler:stream_out_ready
	wire         video_chroma_resampler_avalon_chroma_source_startofpacket;                         // video_chroma_resampler:stream_out_startofpacket -> video_csc:stream_in_startofpacket
	wire         video_chroma_resampler_avalon_chroma_source_endofpacket;                           // video_chroma_resampler:stream_out_endofpacket -> video_csc:stream_in_endofpacket
	wire         video_clipper_normal_avalon_clipper_source_valid;                                  // video_clipper_normal:stream_out_valid -> video_scaler_normal:stream_in_valid
	wire  [15:0] video_clipper_normal_avalon_clipper_source_data;                                   // video_clipper_normal:stream_out_data -> video_scaler_normal:stream_in_data
	wire         video_clipper_normal_avalon_clipper_source_ready;                                  // video_scaler_normal:stream_in_ready -> video_clipper_normal:stream_out_ready
	wire         video_clipper_normal_avalon_clipper_source_startofpacket;                          // video_clipper_normal:stream_out_startofpacket -> video_scaler_normal:stream_in_startofpacket
	wire         video_clipper_normal_avalon_clipper_source_endofpacket;                            // video_clipper_normal:stream_out_endofpacket -> video_scaler_normal:stream_in_endofpacket
	wire         video_csc_avalon_csc_source_valid;                                                 // video_csc:stream_out_valid -> video_rgb_resampler:stream_in_valid
	wire  [23:0] video_csc_avalon_csc_source_data;                                                  // video_csc:stream_out_data -> video_rgb_resampler:stream_in_data
	wire         video_csc_avalon_csc_source_ready;                                                 // video_rgb_resampler:stream_in_ready -> video_csc:stream_out_ready
	wire         video_csc_avalon_csc_source_startofpacket;                                         // video_csc:stream_out_startofpacket -> video_rgb_resampler:stream_in_startofpacket
	wire         video_csc_avalon_csc_source_endofpacket;                                           // video_csc:stream_out_endofpacket -> video_rgb_resampler:stream_in_endofpacket
	wire         mtl_dual_clock_buffer_avalon_dc_buffer_source_valid;                               // mtl_dual_clock_buffer:stream_out_valid -> mtl_controller:valid
	wire  [29:0] mtl_dual_clock_buffer_avalon_dc_buffer_source_data;                                // mtl_dual_clock_buffer:stream_out_data -> mtl_controller:data
	wire         mtl_dual_clock_buffer_avalon_dc_buffer_source_ready;                               // mtl_controller:ready -> mtl_dual_clock_buffer:stream_out_ready
	wire         mtl_dual_clock_buffer_avalon_dc_buffer_source_startofpacket;                       // mtl_dual_clock_buffer:stream_out_startofpacket -> mtl_controller:startofpacket
	wire         mtl_dual_clock_buffer_avalon_dc_buffer_source_endofpacket;                         // mtl_dual_clock_buffer:stream_out_endofpacket -> mtl_controller:endofpacket
	wire         video_decoder_avalon_decoder_source_valid;                                         // video_decoder:stream_out_valid -> video_chroma_resampler:stream_in_valid
	wire  [15:0] video_decoder_avalon_decoder_source_data;                                          // video_decoder:stream_out_data -> video_chroma_resampler:stream_in_data
	wire         video_decoder_avalon_decoder_source_ready;                                         // video_chroma_resampler:stream_in_ready -> video_decoder:stream_out_ready
	wire         video_decoder_avalon_decoder_source_startofpacket;                                 // video_decoder:stream_out_startofpacket -> video_chroma_resampler:stream_in_startofpacket
	wire         video_decoder_avalon_decoder_source_endofpacket;                                   // video_decoder:stream_out_endofpacket -> video_chroma_resampler:stream_in_endofpacket
	wire         pixel_buffer_dma_green_avalon_pixel_source_valid;                                  // pixel_buffer_dma_green:stream_valid -> rgb_resampler_green:stream_in_valid
	wire  [15:0] pixel_buffer_dma_green_avalon_pixel_source_data;                                   // pixel_buffer_dma_green:stream_data -> rgb_resampler_green:stream_in_data
	wire         pixel_buffer_dma_green_avalon_pixel_source_ready;                                  // rgb_resampler_green:stream_in_ready -> pixel_buffer_dma_green:stream_ready
	wire         pixel_buffer_dma_green_avalon_pixel_source_startofpacket;                          // pixel_buffer_dma_green:stream_startofpacket -> rgb_resampler_green:stream_in_startofpacket
	wire         pixel_buffer_dma_green_avalon_pixel_source_endofpacket;                            // pixel_buffer_dma_green:stream_endofpacket -> rgb_resampler_green:stream_in_endofpacket
	wire         video_rgb_resampler_avalon_rgb_source_valid;                                       // video_rgb_resampler:stream_out_valid -> video_clipper_normal:stream_in_valid
	wire  [15:0] video_rgb_resampler_avalon_rgb_source_data;                                        // video_rgb_resampler:stream_out_data -> video_clipper_normal:stream_in_data
	wire         video_rgb_resampler_avalon_rgb_source_ready;                                       // video_clipper_normal:stream_in_ready -> video_rgb_resampler:stream_out_ready
	wire         video_rgb_resampler_avalon_rgb_source_startofpacket;                               // video_rgb_resampler:stream_out_startofpacket -> video_clipper_normal:stream_in_startofpacket
	wire         video_rgb_resampler_avalon_rgb_source_endofpacket;                                 // video_rgb_resampler:stream_out_endofpacket -> video_clipper_normal:stream_in_endofpacket
	wire         rgb_resampler_green_avalon_rgb_source_valid;                                       // rgb_resampler_green:stream_out_valid -> scaler_green:stream_in_valid
	wire  [29:0] rgb_resampler_green_avalon_rgb_source_data;                                        // rgb_resampler_green:stream_out_data -> scaler_green:stream_in_data
	wire         rgb_resampler_green_avalon_rgb_source_ready;                                       // scaler_green:stream_in_ready -> rgb_resampler_green:stream_out_ready
	wire         rgb_resampler_green_avalon_rgb_source_startofpacket;                               // rgb_resampler_green:stream_out_startofpacket -> scaler_green:stream_in_startofpacket
	wire         rgb_resampler_green_avalon_rgb_source_endofpacket;                                 // rgb_resampler_green:stream_out_endofpacket -> scaler_green:stream_in_endofpacket
	wire         video_scaler_normal_avalon_scaler_source_valid;                                    // video_scaler_normal:stream_out_valid -> video_dma_controller_normal:stream_valid
	wire  [15:0] video_scaler_normal_avalon_scaler_source_data;                                     // video_scaler_normal:stream_out_data -> video_dma_controller_normal:stream_data
	wire         video_scaler_normal_avalon_scaler_source_ready;                                    // video_dma_controller_normal:stream_ready -> video_scaler_normal:stream_out_ready
	wire         video_scaler_normal_avalon_scaler_source_startofpacket;                            // video_scaler_normal:stream_out_startofpacket -> video_dma_controller_normal:stream_startofpacket
	wire         video_scaler_normal_avalon_scaler_source_endofpacket;                              // video_scaler_normal:stream_out_endofpacket -> video_dma_controller_normal:stream_endofpacket
	wire         flash_controller_tcm_data_outen;                                                   // flash_controller:tcm_data_outen -> flash_bridge:tcs_tcm_data_outen
	wire         flash_controller_tcm_request;                                                      // flash_controller:tcm_request -> flash_bridge:request
	wire         flash_controller_tcm_write_n_out;                                                  // flash_controller:tcm_write_n_out -> flash_bridge:tcs_tcm_write_n_out
	wire         flash_controller_tcm_read_n_out;                                                   // flash_controller:tcm_read_n_out -> flash_bridge:tcs_tcm_read_n_out
	wire         flash_controller_tcm_grant;                                                        // flash_bridge:grant -> flash_controller:tcm_grant
	wire         flash_controller_tcm_chipselect_n_out;                                             // flash_controller:tcm_chipselect_n_out -> flash_bridge:tcs_tcm_chipselect_n_out
	wire  [22:0] flash_controller_tcm_address_out;                                                  // flash_controller:tcm_address_out -> flash_bridge:tcs_tcm_address_out
	wire   [7:0] flash_controller_tcm_data_out;                                                     // flash_controller:tcm_data_out -> flash_bridge:tcs_tcm_data_out
	wire   [7:0] flash_controller_tcm_data_in;                                                      // flash_bridge:tcs_tcm_data_in -> flash_controller:tcm_data_in
	wire         video_dma_controller_normal_avalon_dma_master_waitrequest;                         // mm_interconnect_0:video_dma_controller_normal_avalon_dma_master_waitrequest -> video_dma_controller_normal:master_waitrequest
	wire  [31:0] video_dma_controller_normal_avalon_dma_master_address;                             // video_dma_controller_normal:master_address -> mm_interconnect_0:video_dma_controller_normal_avalon_dma_master_address
	wire         video_dma_controller_normal_avalon_dma_master_write;                               // video_dma_controller_normal:master_write -> mm_interconnect_0:video_dma_controller_normal_avalon_dma_master_write
	wire  [15:0] video_dma_controller_normal_avalon_dma_master_writedata;                           // video_dma_controller_normal:master_writedata -> mm_interconnect_0:video_dma_controller_normal_avalon_dma_master_writedata
	wire         pixel_buffer_dma_green_avalon_pixel_dma_master_waitrequest;                        // mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_waitrequest -> pixel_buffer_dma_green:master_waitrequest
	wire  [15:0] pixel_buffer_dma_green_avalon_pixel_dma_master_readdata;                           // mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_readdata -> pixel_buffer_dma_green:master_readdata
	wire  [31:0] pixel_buffer_dma_green_avalon_pixel_dma_master_address;                            // pixel_buffer_dma_green:master_address -> mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_address
	wire         pixel_buffer_dma_green_avalon_pixel_dma_master_read;                               // pixel_buffer_dma_green:master_read -> mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_read
	wire         pixel_buffer_dma_green_avalon_pixel_dma_master_readdatavalid;                      // mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_readdatavalid -> pixel_buffer_dma_green:master_readdatavalid
	wire         pixel_buffer_dma_green_avalon_pixel_dma_master_lock;                               // pixel_buffer_dma_green:master_arbiterlock -> mm_interconnect_0:pixel_buffer_dma_green_avalon_pixel_dma_master_lock
	wire  [31:0] cpu_data_master_readdata;                                                          // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                                       // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                                       // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [28:0] cpu_data_master_address;                                                           // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                                        // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                                              // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                                                     // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                                             // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                                         // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                                                   // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                                                // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [27:0] cpu_instruction_master_address;                                                    // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                                       // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                                              // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_readdata;                                 // sram:readdata -> mm_interconnect_0:sram_avalon_sram_slave_readdata
	wire  [19:0] mm_interconnect_0_sram_avalon_sram_slave_address;                                  // mm_interconnect_0:sram_avalon_sram_slave_address -> sram:address
	wire         mm_interconnect_0_sram_avalon_sram_slave_read;                                     // mm_interconnect_0:sram_avalon_sram_slave_read -> sram:read
	wire   [1:0] mm_interconnect_0_sram_avalon_sram_slave_byteenable;                               // mm_interconnect_0:sram_avalon_sram_slave_byteenable -> sram:byteenable
	wire         mm_interconnect_0_sram_avalon_sram_slave_readdatavalid;                            // sram:readdatavalid -> mm_interconnect_0:sram_avalon_sram_slave_readdatavalid
	wire         mm_interconnect_0_sram_avalon_sram_slave_write;                                    // mm_interconnect_0:sram_avalon_sram_slave_write -> sram:write
	wire  [15:0] mm_interconnect_0_sram_avalon_sram_slave_writedata;                                // mm_interconnect_0:sram_avalon_sram_slave_writedata -> sram:writedata
	wire         mm_interconnect_0_audio_avalon_audio_slave_chipselect;                             // mm_interconnect_0:audio_avalon_audio_slave_chipselect -> audio:chipselect
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_readdata;                               // audio:readdata -> mm_interconnect_0:audio_avalon_audio_slave_readdata
	wire   [1:0] mm_interconnect_0_audio_avalon_audio_slave_address;                                // mm_interconnect_0:audio_avalon_audio_slave_address -> audio:address
	wire         mm_interconnect_0_audio_avalon_audio_slave_read;                                   // mm_interconnect_0:audio_avalon_audio_slave_read -> audio:read
	wire         mm_interconnect_0_audio_avalon_audio_slave_write;                                  // mm_interconnect_0:audio_avalon_audio_slave_write -> audio:write
	wire  [31:0] mm_interconnect_0_audio_avalon_audio_slave_writedata;                              // mm_interconnect_0:audio_avalon_audio_slave_writedata -> audio:writedata
	wire  [31:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata;          // audio_and_video_config:readdata -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_readdata
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest;       // audio_and_video_config:waitrequest -> mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_waitrequest
	wire   [1:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address;           // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_address -> audio_and_video_config:address
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read;              // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_read -> audio_and_video_config:read
	wire   [3:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable;        // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_byteenable -> audio_and_video_config:byteenable
	wire         mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write;             // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_write -> audio_and_video_config:write
	wire  [31:0] mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata;         // mm_interconnect_0:audio_and_video_config_avalon_av_config_slave_writedata -> audio_and_video_config:writedata
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_chipselect;             // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_chipselect -> mtl_char_buffer:buf_chipselect
	wire   [7:0] mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_readdata;               // mtl_char_buffer:buf_readdata -> mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_readdata
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_waitrequest;            // mtl_char_buffer:buf_waitrequest -> mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_waitrequest
	wire  [10:0] mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_address;                // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_address -> mtl_char_buffer:buf_address
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_read;                   // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_read -> mtl_char_buffer:buf_read
	wire   [0:0] mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_byteenable;             // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_byteenable -> mtl_char_buffer:buf_byteenable
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_write;                  // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_write -> mtl_char_buffer:buf_write
	wire   [7:0] mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_writedata;              // mm_interconnect_0:mtl_char_buffer_avalon_char_buffer_slave_writedata -> mtl_char_buffer:buf_writedata
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_chipselect;            // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_chipselect -> mtl_char_buffer:ctrl_chipselect
	wire  [31:0] mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_readdata;              // mtl_char_buffer:ctrl_readdata -> mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_readdata
	wire   [0:0] mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_address;               // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_address -> mtl_char_buffer:ctrl_address
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_read;                  // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_read -> mtl_char_buffer:ctrl_read
	wire   [3:0] mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_byteenable;            // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_byteenable -> mtl_char_buffer:ctrl_byteenable
	wire         mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_write;                 // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_write -> mtl_char_buffer:ctrl_write
	wire  [31:0] mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_writedata;             // mm_interconnect_0:mtl_char_buffer_avalon_char_control_slave_writedata -> mtl_char_buffer:ctrl_writedata
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_readdata;            // pixel_buffer_dma_green:slave_readdata -> mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_address;             // mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_address -> pixel_buffer_dma_green:slave_address
	wire         mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_read;                // mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_read -> pixel_buffer_dma_green:slave_read
	wire   [3:0] mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_byteenable;          // mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_byteenable -> pixel_buffer_dma_green:slave_byteenable
	wire         mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_write;               // mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_write -> pixel_buffer_dma_green:slave_write
	wire  [31:0] mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_writedata;           // mm_interconnect_0:pixel_buffer_dma_green_avalon_control_slave_writedata -> pixel_buffer_dma_green:slave_writedata
	wire  [31:0] mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_readdata;   // video_dma_controller_normal:slave_readdata -> mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_address;    // mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_address -> video_dma_controller_normal:slave_address
	wire         mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_read;       // mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_read -> video_dma_controller_normal:slave_read
	wire   [3:0] mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_byteenable; // mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_byteenable -> video_dma_controller_normal:slave_byteenable
	wire         mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_write;      // mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_write -> video_dma_controller_normal:slave_write
	wire  [31:0] mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_writedata;  // mm_interconnect_0:video_dma_controller_normal_avalon_dma_control_slave_writedata -> video_dma_controller_normal:slave_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;                          // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;                            // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;                         // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;                             // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;                                // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;                               // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;                           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_char_lcd_avalon_lcd_slave_chipselect;                            // mm_interconnect_0:char_lcd_avalon_lcd_slave_chipselect -> char_lcd:chipselect
	wire   [7:0] mm_interconnect_0_char_lcd_avalon_lcd_slave_readdata;                              // char_lcd:readdata -> mm_interconnect_0:char_lcd_avalon_lcd_slave_readdata
	wire         mm_interconnect_0_char_lcd_avalon_lcd_slave_waitrequest;                           // char_lcd:waitrequest -> mm_interconnect_0:char_lcd_avalon_lcd_slave_waitrequest
	wire   [0:0] mm_interconnect_0_char_lcd_avalon_lcd_slave_address;                               // mm_interconnect_0:char_lcd_avalon_lcd_slave_address -> char_lcd:address
	wire         mm_interconnect_0_char_lcd_avalon_lcd_slave_read;                                  // mm_interconnect_0:char_lcd_avalon_lcd_slave_read -> char_lcd:read
	wire         mm_interconnect_0_char_lcd_avalon_lcd_slave_write;                                 // mm_interconnect_0:char_lcd_avalon_lcd_slave_write -> char_lcd:write
	wire   [7:0] mm_interconnect_0_char_lcd_avalon_lcd_slave_writedata;                             // mm_interconnect_0:char_lcd_avalon_lcd_slave_writedata -> char_lcd:writedata
	wire         mm_interconnect_0_green_led_avalon_parallel_port_slave_chipselect;                 // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_chipselect -> Green_LED:chipselect
	wire  [31:0] mm_interconnect_0_green_led_avalon_parallel_port_slave_readdata;                   // Green_LED:readdata -> mm_interconnect_0:Green_LED_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_green_led_avalon_parallel_port_slave_address;                    // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_address -> Green_LED:address
	wire         mm_interconnect_0_green_led_avalon_parallel_port_slave_read;                       // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_read -> Green_LED:read
	wire   [3:0] mm_interconnect_0_green_led_avalon_parallel_port_slave_byteenable;                 // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_byteenable -> Green_LED:byteenable
	wire         mm_interconnect_0_green_led_avalon_parallel_port_slave_write;                      // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_write -> Green_LED:write
	wire  [31:0] mm_interconnect_0_green_led_avalon_parallel_port_slave_writedata;                  // mm_interconnect_0:Green_LED_avalon_parallel_port_slave_writedata -> Green_LED:writedata
	wire         mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect;                  // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_chipselect -> red_LEDs:chipselect
	wire  [31:0] mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata;                    // red_LEDs:readdata -> mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_red_leds_avalon_parallel_port_slave_address;                     // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_address -> red_LEDs:address
	wire         mm_interconnect_0_red_leds_avalon_parallel_port_slave_read;                        // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_read -> red_LEDs:read
	wire   [3:0] mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable;                  // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_byteenable -> red_LEDs:byteenable
	wire         mm_interconnect_0_red_leds_avalon_parallel_port_slave_write;                       // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_write -> red_LEDs:write
	wire  [31:0] mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata;                   // mm_interconnect_0:red_LEDs_avalon_parallel_port_slave_writedata -> red_LEDs:writedata
	wire         mm_interconnect_0_switches_avalon_parallel_port_slave_chipselect;                  // mm_interconnect_0:switches_avalon_parallel_port_slave_chipselect -> switches:chipselect
	wire  [31:0] mm_interconnect_0_switches_avalon_parallel_port_slave_readdata;                    // switches:readdata -> mm_interconnect_0:switches_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_switches_avalon_parallel_port_slave_address;                     // mm_interconnect_0:switches_avalon_parallel_port_slave_address -> switches:address
	wire         mm_interconnect_0_switches_avalon_parallel_port_slave_read;                        // mm_interconnect_0:switches_avalon_parallel_port_slave_read -> switches:read
	wire   [3:0] mm_interconnect_0_switches_avalon_parallel_port_slave_byteenable;                  // mm_interconnect_0:switches_avalon_parallel_port_slave_byteenable -> switches:byteenable
	wire         mm_interconnect_0_switches_avalon_parallel_port_slave_write;                       // mm_interconnect_0:switches_avalon_parallel_port_slave_write -> switches:write
	wire  [31:0] mm_interconnect_0_switches_avalon_parallel_port_slave_writedata;                   // mm_interconnect_0:switches_avalon_parallel_port_slave_writedata -> switches:writedata
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect;               // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_chipselect -> pushbuttons:chipselect
	wire  [31:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata;                 // pushbuttons:readdata -> mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address;                  // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_address -> pushbuttons:address
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read;                     // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_read -> pushbuttons:read
	wire   [3:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable;               // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_byteenable -> pushbuttons:byteenable
	wire         mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write;                    // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_write -> pushbuttons:write
	wire  [31:0] mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata;                // mm_interconnect_0:pushbuttons_avalon_parallel_port_slave_writedata -> pushbuttons:writedata
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect;                 // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata;                   // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address;                    // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read;                       // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_read -> HEX3_HEX0:read
	wire   [3:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable;                 // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_byteenable -> HEX3_HEX0:byteenable
	wire         mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write;                      // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_write -> HEX3_HEX0:write
	wire  [31:0] mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata;                  // mm_interconnect_0:HEX3_HEX0_avalon_parallel_port_slave_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_chipselect;                 // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_chipselect -> HEX7_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_readdata;                   // HEX7_HEX4:readdata -> mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_readdata
	wire   [1:0] mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_address;                    // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_address -> HEX7_HEX4:address
	wire         mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_read;                       // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_read -> HEX7_HEX4:read
	wire   [3:0] mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_byteenable;                 // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_byteenable -> HEX7_HEX4:byteenable
	wire         mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_write;                      // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_write -> HEX7_HEX4:write
	wire  [31:0] mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_writedata;                  // mm_interconnect_0:HEX7_HEX4_avalon_parallel_port_slave_writedata -> HEX7_HEX4:writedata
	wire         mm_interconnect_0_ps2_key_avalon_ps2_slave_chipselect;                             // mm_interconnect_0:ps2_key_avalon_ps2_slave_chipselect -> ps2_key:chipselect
	wire  [31:0] mm_interconnect_0_ps2_key_avalon_ps2_slave_readdata;                               // ps2_key:readdata -> mm_interconnect_0:ps2_key_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_key_avalon_ps2_slave_waitrequest;                            // ps2_key:waitrequest -> mm_interconnect_0:ps2_key_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_key_avalon_ps2_slave_address;                                // mm_interconnect_0:ps2_key_avalon_ps2_slave_address -> ps2_key:address
	wire         mm_interconnect_0_ps2_key_avalon_ps2_slave_read;                                   // mm_interconnect_0:ps2_key_avalon_ps2_slave_read -> ps2_key:read
	wire   [3:0] mm_interconnect_0_ps2_key_avalon_ps2_slave_byteenable;                             // mm_interconnect_0:ps2_key_avalon_ps2_slave_byteenable -> ps2_key:byteenable
	wire         mm_interconnect_0_ps2_key_avalon_ps2_slave_write;                                  // mm_interconnect_0:ps2_key_avalon_ps2_slave_write -> ps2_key:write
	wire  [31:0] mm_interconnect_0_ps2_key_avalon_ps2_slave_writedata;                              // mm_interconnect_0:ps2_key_avalon_ps2_slave_writedata -> ps2_key:writedata
	wire         mm_interconnect_0_ps2_mouse_avalon_ps2_slave_chipselect;                           // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_chipselect -> ps2_mouse:chipselect
	wire  [31:0] mm_interconnect_0_ps2_mouse_avalon_ps2_slave_readdata;                             // ps2_mouse:readdata -> mm_interconnect_0:ps2_mouse_avalon_ps2_slave_readdata
	wire         mm_interconnect_0_ps2_mouse_avalon_ps2_slave_waitrequest;                          // ps2_mouse:waitrequest -> mm_interconnect_0:ps2_mouse_avalon_ps2_slave_waitrequest
	wire   [0:0] mm_interconnect_0_ps2_mouse_avalon_ps2_slave_address;                              // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_address -> ps2_mouse:address
	wire         mm_interconnect_0_ps2_mouse_avalon_ps2_slave_read;                                 // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_read -> ps2_mouse:read
	wire   [3:0] mm_interconnect_0_ps2_mouse_avalon_ps2_slave_byteenable;                           // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_byteenable -> ps2_mouse:byteenable
	wire         mm_interconnect_0_ps2_mouse_avalon_ps2_slave_write;                                // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_write -> ps2_mouse:write
	wire  [31:0] mm_interconnect_0_ps2_mouse_avalon_ps2_slave_writedata;                            // mm_interconnect_0:ps2_mouse_avalon_ps2_slave_writedata -> ps2_mouse:writedata
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect;                       // mm_interconnect_0:serial_port_avalon_rs232_slave_chipselect -> serial_port:chipselect
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_readdata;                         // serial_port:readdata -> mm_interconnect_0:serial_port_avalon_rs232_slave_readdata
	wire   [0:0] mm_interconnect_0_serial_port_avalon_rs232_slave_address;                          // mm_interconnect_0:serial_port_avalon_rs232_slave_address -> serial_port:address
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_read;                             // mm_interconnect_0:serial_port_avalon_rs232_slave_read -> serial_port:read
	wire   [3:0] mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable;                       // mm_interconnect_0:serial_port_avalon_rs232_slave_byteenable -> serial_port:byteenable
	wire         mm_interconnect_0_serial_port_avalon_rs232_slave_write;                            // mm_interconnect_0:serial_port_avalon_rs232_slave_write -> serial_port:write
	wire  [31:0] mm_interconnect_0_serial_port_avalon_rs232_slave_writedata;                        // mm_interconnect_0:serial_port_avalon_rs232_slave_writedata -> serial_port:writedata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect;                          // mm_interconnect_0:sd_card_avalon_sdcard_slave_chipselect -> sd_card:i_avalon_chip_select
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata;                            // sd_card:o_avalon_readdata -> mm_interconnect_0:sd_card_avalon_sdcard_slave_readdata
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest;                         // sd_card:o_avalon_waitrequest -> mm_interconnect_0:sd_card_avalon_sdcard_slave_waitrequest
	wire   [7:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_address;                             // mm_interconnect_0:sd_card_avalon_sdcard_slave_address -> sd_card:i_avalon_address
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_read;                                // mm_interconnect_0:sd_card_avalon_sdcard_slave_read -> sd_card:i_avalon_read
	wire   [3:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable;                          // mm_interconnect_0:sd_card_avalon_sdcard_slave_byteenable -> sd_card:i_avalon_byteenable
	wire         mm_interconnect_0_sd_card_avalon_sdcard_slave_write;                               // mm_interconnect_0:sd_card_avalon_sdcard_slave_write -> sd_card:i_avalon_write
	wire  [31:0] mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata;                           // mm_interconnect_0:sd_card_avalon_sdcard_slave_writedata -> sd_card:i_avalon_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                                    // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                                     // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_readdata;                      // performance_counter:readdata -> mm_interconnect_0:performance_counter_control_slave_readdata
	wire   [3:0] mm_interconnect_0_performance_counter_control_slave_address;                       // mm_interconnect_0:performance_counter_control_slave_address -> performance_counter:address
	wire         mm_interconnect_0_performance_counter_control_slave_begintransfer;                 // mm_interconnect_0:performance_counter_control_slave_begintransfer -> performance_counter:begintransfer
	wire         mm_interconnect_0_performance_counter_control_slave_write;                         // mm_interconnect_0:performance_counter_control_slave_write -> performance_counter:write
	wire  [31:0] mm_interconnect_0_performance_counter_control_slave_writedata;                     // mm_interconnect_0:performance_counter_control_slave_writedata -> performance_counter:writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;                                    // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;                                 // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;                                 // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;                                     // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                                        // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;                                  // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;                                       // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;                                   // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                                             // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                                               // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                            // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                                                // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                                                   // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                                             // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                          // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                                                  // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                                              // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_onchip_memory_s1_chipselect;                                     // mm_interconnect_0:onchip_memory_s1_chipselect -> onchip_memory:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_readdata;                                       // onchip_memory:readdata -> mm_interconnect_0:onchip_memory_s1_readdata
	wire  [12:0] mm_interconnect_0_onchip_memory_s1_address;                                        // mm_interconnect_0:onchip_memory_s1_address -> onchip_memory:address
	wire   [3:0] mm_interconnect_0_onchip_memory_s1_byteenable;                                     // mm_interconnect_0:onchip_memory_s1_byteenable -> onchip_memory:byteenable
	wire         mm_interconnect_0_onchip_memory_s1_write;                                          // mm_interconnect_0:onchip_memory_s1_write -> onchip_memory:write
	wire  [31:0] mm_interconnect_0_onchip_memory_s1_writedata;                                      // mm_interconnect_0:onchip_memory_s1_writedata -> onchip_memory:writedata
	wire         mm_interconnect_0_onchip_memory_s1_clken;                                          // mm_interconnect_0:onchip_memory_s1_clken -> onchip_memory:clken
	wire         mm_interconnect_0_timer_s1_chipselect;                                             // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                                               // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                                                // mm_interconnect_0:timer_s1_address -> timer:address
	wire         mm_interconnect_0_timer_s1_write;                                                  // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                                              // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire   [7:0] mm_interconnect_0_flash_controller_uas_readdata;                                   // flash_controller:uas_readdata -> mm_interconnect_0:flash_controller_uas_readdata
	wire         mm_interconnect_0_flash_controller_uas_waitrequest;                                // flash_controller:uas_waitrequest -> mm_interconnect_0:flash_controller_uas_waitrequest
	wire         mm_interconnect_0_flash_controller_uas_debugaccess;                                // mm_interconnect_0:flash_controller_uas_debugaccess -> flash_controller:uas_debugaccess
	wire  [22:0] mm_interconnect_0_flash_controller_uas_address;                                    // mm_interconnect_0:flash_controller_uas_address -> flash_controller:uas_address
	wire         mm_interconnect_0_flash_controller_uas_read;                                       // mm_interconnect_0:flash_controller_uas_read -> flash_controller:uas_read
	wire   [0:0] mm_interconnect_0_flash_controller_uas_byteenable;                                 // mm_interconnect_0:flash_controller_uas_byteenable -> flash_controller:uas_byteenable
	wire         mm_interconnect_0_flash_controller_uas_readdatavalid;                              // flash_controller:uas_readdatavalid -> mm_interconnect_0:flash_controller_uas_readdatavalid
	wire         mm_interconnect_0_flash_controller_uas_lock;                                       // mm_interconnect_0:flash_controller_uas_lock -> flash_controller:uas_lock
	wire         mm_interconnect_0_flash_controller_uas_write;                                      // mm_interconnect_0:flash_controller_uas_write -> flash_controller:uas_write
	wire   [7:0] mm_interconnect_0_flash_controller_uas_writedata;                                  // mm_interconnect_0:flash_controller_uas_writedata -> flash_controller:uas_writedata
	wire   [0:0] mm_interconnect_0_flash_controller_uas_burstcount;                                 // mm_interconnect_0:flash_controller_uas_burstcount -> flash_controller:uas_burstcount
	wire         irq_mapper_receiver0_irq;                                                          // pushbuttons:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                          // switches:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                          // audio:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                          // ps2_key:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                          // ps2_mouse:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                          // serial_port:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                          // jtag_uart:av_irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                                          // timer:irq -> irq_mapper:receiver7_irq
	wire  [31:0] cpu_irq_irq;                                                                       // irq_mapper:sender_irq -> cpu:irq
	wire         scaler_green_avalon_scaler_source_valid;                                           // scaler_green:stream_out_valid -> avalon_st_adapter:in_0_valid
	wire  [29:0] scaler_green_avalon_scaler_source_data;                                            // scaler_green:stream_out_data -> avalon_st_adapter:in_0_data
	wire         scaler_green_avalon_scaler_source_ready;                                           // avalon_st_adapter:in_0_ready -> scaler_green:stream_out_ready
	wire   [1:0] scaler_green_avalon_scaler_source_channel;                                         // scaler_green:stream_out_channel -> avalon_st_adapter:in_0_channel
	wire         scaler_green_avalon_scaler_source_startofpacket;                                   // scaler_green:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	wire         scaler_green_avalon_scaler_source_endofpacket;                                     // scaler_green:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	wire         avalon_st_adapter_out_0_valid;                                                     // avalon_st_adapter:out_0_valid -> alpha_blending:background_valid
	wire  [29:0] avalon_st_adapter_out_0_data;                                                      // avalon_st_adapter:out_0_data -> alpha_blending:background_data
	wire         avalon_st_adapter_out_0_ready;                                                     // alpha_blending:background_ready -> avalon_st_adapter:out_0_ready
	wire         avalon_st_adapter_out_0_startofpacket;                                             // avalon_st_adapter:out_0_startofpacket -> alpha_blending:background_startofpacket
	wire         avalon_st_adapter_out_0_endofpacket;                                               // avalon_st_adapter:out_0_endofpacket -> alpha_blending:background_endofpacket
	wire         rst_controller_reset_out_reset;                                                    // rst_controller:reset_out -> [Green_LED:reset, HEX3_HEX0:reset, HEX7_HEX4:reset, alpha_blending:reset, audio:reset, audio_and_video_config:reset, avalon_st_adapter:in_rst_0_reset, char_lcd:reset, cpu:reset_n, flash_bridge:reset, flash_controller:reset_reset, irq_mapper:reset, jtag_uart:rst_n, mm_interconnect_0:video_dma_controller_normal_reset_reset_bridge_in_reset_reset, mtl_char_buffer:reset, mtl_dual_clock_buffer:reset_stream_in, onchip_memory:reset, performance_counter:reset_n, pixel_buffer_dma_green:reset, ps2_key:reset, ps2_mouse:reset, pushbuttons:reset, red_LEDs:reset, rgb_resampler_green:reset, rst_translator:in_reset, scaler_green:reset, sd_card:i_reset_n, sdram:reset_n, serial_port:reset, sram:reset, switches:reset, sysid:reset_n, timer:reset_n, video_chroma_resampler:reset, video_clipper_normal:reset, video_csc:reset, video_decoder:reset, video_dma_controller_normal:reset, video_rgb_resampler:reset, video_scaler_normal:reset]
	wire         rst_controller_reset_out_reset_req;                                                // rst_controller:reset_req -> [cpu:reset_req, onchip_memory:reset_req, rst_translator:reset_req_in]
	wire         cpu_debug_reset_request_reset;                                                     // cpu:debug_reset_request -> [rst_controller:reset_in0, rst_controller_002:reset_in0]
	wire         sys_sdram_pll_reset_source_reset;                                                  // sys_sdram_pll:reset_source_reset -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                                                // rst_controller_001:reset_out -> audio_pll:ref_reset_reset
	wire         rst_controller_002_reset_out_reset;                                                // rst_controller_002:reset_out -> [mtl_controller:reset, mtl_dual_clock_buffer:reset_stream_out]
	wire         video_pll_reset_source_reset;                                                      // video_pll:reset_source_reset -> rst_controller_002:reset_in1
	wire         rst_controller_003_reset_out_reset;                                                // rst_controller_003:reset_out -> sys_sdram_pll:ref_reset_reset
	wire         rst_controller_004_reset_out_reset;                                                // rst_controller_004:reset_out -> video_pll:ref_reset_reset

	nios_system_Green_LED green_led (
		.clk        (sys_clk_out_clk),                                                   //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                    //                      reset.reset
		.address    (mm_interconnect_0_green_led_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_green_led_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_green_led_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_green_led_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_green_led_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_green_led_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_green_led_avalon_parallel_port_slave_readdata),   //                           .readdata
		.LEDG       (green_led_external_interface_export)                                //         external_interface.export
	);

	nios_system_HEX3_HEX0 hex3_hex0 (
		.clk        (sys_clk_out_clk),                                                   //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                    //                      reset.reset
		.address    (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata),   //                           .readdata
		.HEX0       (hex3_hex0_external_interface_HEX0),                                 //         external_interface.export
		.HEX1       (hex3_hex0_external_interface_HEX1),                                 //                           .export
		.HEX2       (hex3_hex0_external_interface_HEX2),                                 //                           .export
		.HEX3       (hex3_hex0_external_interface_HEX3)                                  //                           .export
	);

	nios_system_HEX7_HEX4 hex7_hex4 (
		.clk        (sys_clk_out_clk),                                                   //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                    //                      reset.reset
		.address    (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_readdata),   //                           .readdata
		.HEX4       (hex7_hex4_external_interface_HEX4),                                 //         external_interface.export
		.HEX5       (hex7_hex4_external_interface_HEX5),                                 //                           .export
		.HEX6       (hex7_hex4_external_interface_HEX6),                                 //                           .export
		.HEX7       (hex7_hex4_external_interface_HEX7)                                  //                           .export
	);

	nios_system_alpha_blending alpha_blending (
		.clk                      (sys_clk_out_clk),                                    //                    clk.clk
		.reset                    (rst_controller_reset_out_reset),                     //                  reset.reset
		.foreground_data          (mtl_char_buffer_avalon_char_source_data),            // avalon_foreground_sink.data
		.foreground_startofpacket (mtl_char_buffer_avalon_char_source_startofpacket),   //                       .startofpacket
		.foreground_endofpacket   (mtl_char_buffer_avalon_char_source_endofpacket),     //                       .endofpacket
		.foreground_valid         (mtl_char_buffer_avalon_char_source_valid),           //                       .valid
		.foreground_ready         (mtl_char_buffer_avalon_char_source_ready),           //                       .ready
		.background_data          (avalon_st_adapter_out_0_data),                       // avalon_background_sink.data
		.background_startofpacket (avalon_st_adapter_out_0_startofpacket),              //                       .startofpacket
		.background_endofpacket   (avalon_st_adapter_out_0_endofpacket),                //                       .endofpacket
		.background_valid         (avalon_st_adapter_out_0_valid),                      //                       .valid
		.background_ready         (avalon_st_adapter_out_0_ready),                      //                       .ready
		.output_ready             (alpha_blending_avalon_blended_source_ready),         //  avalon_blended_source.ready
		.output_data              (alpha_blending_avalon_blended_source_data),          //                       .data
		.output_startofpacket     (alpha_blending_avalon_blended_source_startofpacket), //                       .startofpacket
		.output_endofpacket       (alpha_blending_avalon_blended_source_endofpacket),   //                       .endofpacket
		.output_valid             (alpha_blending_avalon_blended_source_valid)          //                       .valid
	);

	nios_system_audio audio (
		.clk         (sys_clk_out_clk),                                       //                clk.clk
		.reset       (rst_controller_reset_out_reset),                        //              reset.reset
		.address     (mm_interconnect_0_audio_avalon_audio_slave_address),    // avalon_audio_slave.address
		.chipselect  (mm_interconnect_0_audio_avalon_audio_slave_chipselect), //                   .chipselect
		.read        (mm_interconnect_0_audio_avalon_audio_slave_read),       //                   .read
		.write       (mm_interconnect_0_audio_avalon_audio_slave_write),      //                   .write
		.writedata   (mm_interconnect_0_audio_avalon_audio_slave_writedata),  //                   .writedata
		.readdata    (mm_interconnect_0_audio_avalon_audio_slave_readdata),   //                   .readdata
		.irq         (irq_mapper_receiver2_irq),                              //          interrupt.irq
		.AUD_ADCDAT  (audio_external_interface_ADCDAT),                       // external_interface.export
		.AUD_ADCLRCK (audio_external_interface_ADCLRCK),                      //                   .export
		.AUD_BCLK    (audio_external_interface_BCLK),                         //                   .export
		.AUD_DACDAT  (audio_external_interface_DACDAT),                       //                   .export
		.AUD_DACLRCK (audio_external_interface_DACLRCK)                       //                   .export
	);

	nios_system_audio_and_video_config audio_and_video_config (
		.clk         (sys_clk_out_clk),                                                             //                    clk.clk
		.reset       (rst_controller_reset_out_reset),                                              //                  reset.reset
		.address     (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address),     // avalon_av_config_slave.address
		.byteenable  (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable),  //                       .byteenable
		.read        (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read),        //                       .read
		.write       (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write),       //                       .write
		.writedata   (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata),   //                       .writedata
		.readdata    (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata),    //                       .readdata
		.waitrequest (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest), //                       .waitrequest
		.I2C_SDAT    (audio_and_video_config_external_interface_SDAT),                              //     external_interface.export
		.I2C_SCLK    (audio_and_video_config_external_interface_SCLK)                               //                       .export
	);

	nios_system_audio_pll audio_pll (
		.ref_clk_clk        (clk_50_3_in_clk),                    //      ref_clk.clk
		.ref_reset_reset    (rst_controller_001_reset_out_reset), //    ref_reset.reset
		.audio_clk_clk      (audio_clk_out_clk),                  //    audio_clk.clk
		.reset_source_reset ()                                    // reset_source.reset
	);

	nios_system_char_lcd char_lcd (
		.clk         (sys_clk_out_clk),                                         //                clk.clk
		.reset       (rst_controller_reset_out_reset),                          //              reset.reset
		.address     (mm_interconnect_0_char_lcd_avalon_lcd_slave_address),     //   avalon_lcd_slave.address
		.chipselect  (mm_interconnect_0_char_lcd_avalon_lcd_slave_chipselect),  //                   .chipselect
		.read        (mm_interconnect_0_char_lcd_avalon_lcd_slave_read),        //                   .read
		.write       (mm_interconnect_0_char_lcd_avalon_lcd_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_char_lcd_avalon_lcd_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_char_lcd_avalon_lcd_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_char_lcd_avalon_lcd_slave_waitrequest), //                   .waitrequest
		.LCD_DATA    (char_lcd_external_interface_DATA),                        // external_interface.export
		.LCD_ON      (char_lcd_external_interface_ON),                          //                   .export
		.LCD_BLON    (char_lcd_external_interface_BLON),                        //                   .export
		.LCD_EN      (char_lcd_external_interface_EN),                          //                   .export
		.LCD_RS      (char_lcd_external_interface_RS),                          //                   .export
		.LCD_RW      (char_lcd_external_interface_RW)                           //                   .export
	);

	nios_system_cpu cpu (
		.clk                                 (sys_clk_out_clk),                                   //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                   //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios_system_flash_bridge flash_bridge (
		.clk                      (sys_clk_out_clk),                       //   clk.clk
		.reset                    (rst_controller_reset_out_reset),        // reset.reset
		.request                  (flash_controller_tcm_request),          //   tcs.request
		.grant                    (flash_controller_tcm_grant),            //      .grant
		.tcs_tcm_address_out      (flash_controller_tcm_address_out),      //      .address_out
		.tcs_tcm_read_n_out       (flash_controller_tcm_read_n_out),       //      .read_n_out
		.tcs_tcm_write_n_out      (flash_controller_tcm_write_n_out),      //      .write_n_out
		.tcs_tcm_data_out         (flash_controller_tcm_data_out),         //      .data_out
		.tcs_tcm_data_outen       (flash_controller_tcm_data_outen),       //      .data_outen
		.tcs_tcm_data_in          (flash_controller_tcm_data_in),          //      .data_in
		.tcs_tcm_chipselect_n_out (flash_controller_tcm_chipselect_n_out), //      .chipselect_n_out
		.tcm_address_out          (flash_bridge_out_tcm_address_out),      //   out.tcm_address_out
		.tcm_read_n_out           (flash_bridge_out_tcm_read_n_out),       //      .tcm_read_n_out
		.tcm_write_n_out          (flash_bridge_out_tcm_write_n_out),      //      .tcm_write_n_out
		.tcm_data_out             (flash_bridge_out_tcm_data_out),         //      .tcm_data_out
		.tcm_chipselect_n_out     (flash_bridge_out_tcm_chipselect_n_out)  //      .tcm_chipselect_n_out
	);

	nios_system_flash_controller #(
		.TCM_ADDRESS_W                  (23),
		.TCM_DATA_W                     (8),
		.TCM_BYTEENABLE_W               (1),
		.TCM_READ_WAIT                  (160),
		.TCM_WRITE_WAIT                 (160),
		.TCM_SETUP_WAIT                 (60),
		.TCM_DATA_HOLD                  (60),
		.TCM_TURNAROUND_TIME            (2),
		.TCM_TIMING_UNITS               (0),
		.TCM_READLATENCY                (2),
		.TCM_SYMBOLS_PER_WORD           (1),
		.USE_READDATA                   (1),
		.USE_WRITEDATA                  (1),
		.USE_READ                       (1),
		.USE_WRITE                      (1),
		.USE_BYTEENABLE                 (0),
		.USE_CHIPSELECT                 (1),
		.USE_LOCK                       (0),
		.USE_ADDRESS                    (1),
		.USE_WAITREQUEST                (0),
		.USE_WRITEBYTEENABLE            (0),
		.USE_OUTPUTENABLE               (0),
		.USE_RESETREQUEST               (0),
		.USE_IRQ                        (0),
		.USE_RESET_OUTPUT               (0),
		.ACTIVE_LOW_READ                (1),
		.ACTIVE_LOW_LOCK                (0),
		.ACTIVE_LOW_WRITE               (1),
		.ACTIVE_LOW_CHIPSELECT          (1),
		.ACTIVE_LOW_BYTEENABLE          (0),
		.ACTIVE_LOW_OUTPUTENABLE        (0),
		.ACTIVE_LOW_WRITEBYTEENABLE     (0),
		.ACTIVE_LOW_WAITREQUEST         (0),
		.ACTIVE_LOW_BEGINTRANSFER       (0),
		.CHIPSELECT_THROUGH_READLATENCY (0)
	) flash_controller (
		.clk_clk              (sys_clk_out_clk),                                      //   clk.clk
		.reset_reset          (rst_controller_reset_out_reset),                       // reset.reset
		.uas_address          (mm_interconnect_0_flash_controller_uas_address),       //   uas.address
		.uas_burstcount       (mm_interconnect_0_flash_controller_uas_burstcount),    //      .burstcount
		.uas_read             (mm_interconnect_0_flash_controller_uas_read),          //      .read
		.uas_write            (mm_interconnect_0_flash_controller_uas_write),         //      .write
		.uas_waitrequest      (mm_interconnect_0_flash_controller_uas_waitrequest),   //      .waitrequest
		.uas_readdatavalid    (mm_interconnect_0_flash_controller_uas_readdatavalid), //      .readdatavalid
		.uas_byteenable       (mm_interconnect_0_flash_controller_uas_byteenable),    //      .byteenable
		.uas_readdata         (mm_interconnect_0_flash_controller_uas_readdata),      //      .readdata
		.uas_writedata        (mm_interconnect_0_flash_controller_uas_writedata),     //      .writedata
		.uas_lock             (mm_interconnect_0_flash_controller_uas_lock),          //      .lock
		.uas_debugaccess      (mm_interconnect_0_flash_controller_uas_debugaccess),   //      .debugaccess
		.tcm_write_n_out      (flash_controller_tcm_write_n_out),                     //   tcm.write_n_out
		.tcm_read_n_out       (flash_controller_tcm_read_n_out),                      //      .read_n_out
		.tcm_chipselect_n_out (flash_controller_tcm_chipselect_n_out),                //      .chipselect_n_out
		.tcm_request          (flash_controller_tcm_request),                         //      .request
		.tcm_grant            (flash_controller_tcm_grant),                           //      .grant
		.tcm_address_out      (flash_controller_tcm_address_out),                     //      .address_out
		.tcm_data_out         (flash_controller_tcm_data_out),                        //      .data_out
		.tcm_data_outen       (flash_controller_tcm_data_outen),                      //      .data_outen
		.tcm_data_in          (flash_controller_tcm_data_in)                          //      .data_in
	);

	nios_system_jtag_uart jtag_uart (
		.clk            (sys_clk_out_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver6_irq)                                   //               irq.irq
	);

	nios_system_mtl_char_buffer mtl_char_buffer (
		.clk                  (sys_clk_out_clk),                                                        //                       clk.clk
		.reset                (rst_controller_reset_out_reset),                                         //                     reset.reset
		.ctrl_address         (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_address),    // avalon_char_control_slave.address
		.ctrl_byteenable      (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_byteenable), //                          .byteenable
		.ctrl_chipselect      (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_chipselect), //                          .chipselect
		.ctrl_read            (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_read),       //                          .read
		.ctrl_write           (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_write),      //                          .write
		.ctrl_writedata       (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_writedata),  //                          .writedata
		.ctrl_readdata        (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_readdata),   //                          .readdata
		.buf_byteenable       (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_byteenable),  //  avalon_char_buffer_slave.byteenable
		.buf_chipselect       (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_chipselect),  //                          .chipselect
		.buf_read             (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_read),        //                          .read
		.buf_write            (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_write),       //                          .write
		.buf_writedata        (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_writedata),   //                          .writedata
		.buf_readdata         (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_readdata),    //                          .readdata
		.buf_waitrequest      (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_waitrequest), //                          .waitrequest
		.buf_address          (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_address),     //                          .address
		.stream_ready         (mtl_char_buffer_avalon_char_source_ready),                               //        avalon_char_source.ready
		.stream_startofpacket (mtl_char_buffer_avalon_char_source_startofpacket),                       //                          .startofpacket
		.stream_endofpacket   (mtl_char_buffer_avalon_char_source_endofpacket),                         //                          .endofpacket
		.stream_valid         (mtl_char_buffer_avalon_char_source_valid),                               //                          .valid
		.stream_data          (mtl_char_buffer_avalon_char_source_data)                                 //                          .data
	);

	nios_system_mtl_controller mtl_controller (
		.clk           (mtl_clk_out_clk),                                             //                clk.clk
		.reset         (rst_controller_002_reset_out_reset),                          //              reset.reset
		.data          (mtl_dual_clock_buffer_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (mtl_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (mtl_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (mtl_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (mtl_dual_clock_buffer_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (mtl_controller_external_interface_CLK),                       // external_interface.export
		.VGA_HS        (mtl_controller_external_interface_HS),                        //                   .export
		.VGA_VS        (mtl_controller_external_interface_VS),                        //                   .export
		.VGA_DATA_EN   (mtl_controller_external_interface_DATA_EN),                   //                   .export
		.VGA_R         (mtl_controller_external_interface_R),                         //                   .export
		.VGA_G         (mtl_controller_external_interface_G),                         //                   .export
		.VGA_B         (mtl_controller_external_interface_B)                          //                   .export
	);

	nios_system_mtl_dual_clock_buffer mtl_dual_clock_buffer (
		.clk_stream_in            (sys_clk_out_clk),                                             //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                              //         reset_stream_in.reset
		.clk_stream_out           (mtl_clk_out_clk),                                             //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_002_reset_out_reset),                          //        reset_stream_out.reset
		.stream_in_ready          (alpha_blending_avalon_blended_source_ready),                  //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (alpha_blending_avalon_blended_source_startofpacket),          //                        .startofpacket
		.stream_in_endofpacket    (alpha_blending_avalon_blended_source_endofpacket),            //                        .endofpacket
		.stream_in_valid          (alpha_blending_avalon_blended_source_valid),                  //                        .valid
		.stream_in_data           (alpha_blending_avalon_blended_source_data),                   //                        .data
		.stream_out_ready         (mtl_dual_clock_buffer_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (mtl_dual_clock_buffer_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (mtl_dual_clock_buffer_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (mtl_dual_clock_buffer_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (mtl_dual_clock_buffer_avalon_dc_buffer_source_data)           //                        .data
	);

	nios_system_onchip_memory onchip_memory (
		.clk        (sys_clk_out_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),            //       .reset_req
		.freeze     (1'b0)                                           // (terminated)
	);

	nios_system_performance_counter performance_counter (
		.clk           (sys_clk_out_clk),                                                   //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                   //         reset.reset_n
		.address       (mm_interconnect_0_performance_counter_control_slave_address),       // control_slave.address
		.begintransfer (mm_interconnect_0_performance_counter_control_slave_begintransfer), //              .begintransfer
		.readdata      (mm_interconnect_0_performance_counter_control_slave_readdata),      //              .readdata
		.write         (mm_interconnect_0_performance_counter_control_slave_write),         //              .write
		.writedata     (mm_interconnect_0_performance_counter_control_slave_writedata)      //              .writedata
	);

	nios_system_pixel_buffer_dma_green pixel_buffer_dma_green (
		.clk                  (sys_clk_out_clk),                                                          //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                           //                   reset.reset
		.master_readdatavalid (pixel_buffer_dma_green_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (pixel_buffer_dma_green_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (pixel_buffer_dma_green_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (pixel_buffer_dma_green_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (pixel_buffer_dma_green_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (pixel_buffer_dma_green_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (pixel_buffer_dma_green_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (pixel_buffer_dma_green_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (pixel_buffer_dma_green_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (pixel_buffer_dma_green_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (pixel_buffer_dma_green_avalon_pixel_source_data)                           //                        .data
	);

	nios_system_ps2_key ps2_key (
		.clk         (sys_clk_out_clk),                                        //                clk.clk
		.reset       (rst_controller_reset_out_reset),                         //              reset.reset
		.address     (mm_interconnect_0_ps2_key_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_key_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_key_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_key_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_key_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_key_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_key_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_key_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver3_irq),                               //          interrupt.irq
		.PS2_CLK     (ps2_key_external_interface_CLK),                         // external_interface.export
		.PS2_DAT     (ps2_key_external_interface_DAT)                          //                   .export
	);

	nios_system_ps2_key ps2_mouse (
		.clk         (sys_clk_out_clk),                                          //                clk.clk
		.reset       (rst_controller_reset_out_reset),                           //              reset.reset
		.address     (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_address),     //   avalon_ps2_slave.address
		.chipselect  (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_chipselect),  //                   .chipselect
		.byteenable  (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_byteenable),  //                   .byteenable
		.read        (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_read),        //                   .read
		.write       (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_write),       //                   .write
		.writedata   (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_writedata),   //                   .writedata
		.readdata    (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_readdata),    //                   .readdata
		.waitrequest (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_waitrequest), //                   .waitrequest
		.irq         (irq_mapper_receiver4_irq),                                 //          interrupt.irq
		.PS2_CLK     (ps2_mouse_external_interface_CLK),                         // external_interface.export
		.PS2_DAT     (ps2_mouse_external_interface_DAT)                          //                   .export
	);

	nios_system_pushbuttons pushbuttons (
		.clk        (sys_clk_out_clk),                                                     //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                      //                      reset.reset
		.address    (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata),   //                           .readdata
		.KEY        (pushbuttons_external_interface_export),                               //         external_interface.export
		.irq        (irq_mapper_receiver0_irq)                                             //                  interrupt.irq
	);

	nios_system_red_LEDs red_leds (
		.clk        (sys_clk_out_clk),                                                  //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                   //                      reset.reset
		.address    (mm_interconnect_0_red_leds_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_red_leds_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_red_leds_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata),   //                           .readdata
		.LEDR       (red_leds_external_interface_export)                                //         external_interface.export
	);

	nios_system_rgb_resampler_green rgb_resampler_green (
		.clk                      (sys_clk_out_clk),                                          //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                           //             reset.reset
		.stream_in_startofpacket  (pixel_buffer_dma_green_avalon_pixel_source_startofpacket), //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (pixel_buffer_dma_green_avalon_pixel_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (pixel_buffer_dma_green_avalon_pixel_source_valid),         //                  .valid
		.stream_in_ready          (pixel_buffer_dma_green_avalon_pixel_source_ready),         //                  .ready
		.stream_in_data           (pixel_buffer_dma_green_avalon_pixel_source_data),          //                  .data
		.stream_out_ready         (rgb_resampler_green_avalon_rgb_source_ready),              // avalon_rgb_source.ready
		.stream_out_startofpacket (rgb_resampler_green_avalon_rgb_source_startofpacket),      //                  .startofpacket
		.stream_out_endofpacket   (rgb_resampler_green_avalon_rgb_source_endofpacket),        //                  .endofpacket
		.stream_out_valid         (rgb_resampler_green_avalon_rgb_source_valid),              //                  .valid
		.stream_out_data          (rgb_resampler_green_avalon_rgb_source_data)                //                  .data
	);

	nios_system_scaler_green scaler_green (
		.clk                      (sys_clk_out_clk),                                     //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //                reset.reset
		.stream_in_startofpacket  (rgb_resampler_green_avalon_rgb_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (rgb_resampler_green_avalon_rgb_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (rgb_resampler_green_avalon_rgb_source_valid),         //                     .valid
		.stream_in_ready          (rgb_resampler_green_avalon_rgb_source_ready),         //                     .ready
		.stream_in_data           (rgb_resampler_green_avalon_rgb_source_data),          //                     .data
		.stream_out_ready         (scaler_green_avalon_scaler_source_ready),             // avalon_scaler_source.ready
		.stream_out_startofpacket (scaler_green_avalon_scaler_source_startofpacket),     //                     .startofpacket
		.stream_out_endofpacket   (scaler_green_avalon_scaler_source_endofpacket),       //                     .endofpacket
		.stream_out_valid         (scaler_green_avalon_scaler_source_valid),             //                     .valid
		.stream_out_data          (scaler_green_avalon_scaler_source_data),              //                     .data
		.stream_out_channel       (scaler_green_avalon_scaler_source_channel)            //                     .channel
	);

	Altera_UP_SD_Card_Avalon_Interface sd_card (
		.i_avalon_chip_select (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),  // avalon_sdcard_slave.chipselect
		.i_avalon_address     (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),     //                    .address
		.i_avalon_read        (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),        //                    .read
		.i_avalon_write       (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),       //                    .write
		.i_avalon_byteenable  (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),  //                    .byteenable
		.i_avalon_writedata   (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),   //                    .writedata
		.o_avalon_readdata    (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),    //                    .readdata
		.o_avalon_waitrequest (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest), //                    .waitrequest
		.i_clock              (sys_clk_out_clk),                                           //                 clk.clk
		.i_reset_n            (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.b_SD_cmd             (sd_card_conduit_end_b_SD_cmd),                              //         conduit_end.export
		.b_SD_dat             (sd_card_conduit_end_b_SD_dat),                              //                    .export
		.b_SD_dat3            (sd_card_conduit_end_b_SD_dat3),                             //                    .export
		.o_SD_clock           (sd_card_conduit_end_o_SD_clock)                             //                    .export
	);

	nios_system_sdram sdram (
		.clk            (sys_clk_out_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	nios_system_serial_port serial_port (
		.clk        (sys_clk_out_clk),                                             //                clk.clk
		.reset      (rst_controller_reset_out_reset),                              //              reset.reset
		.address    (mm_interconnect_0_serial_port_avalon_rs232_slave_address),    // avalon_rs232_slave.address
		.chipselect (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect), //                   .chipselect
		.byteenable (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable), //                   .byteenable
		.read       (mm_interconnect_0_serial_port_avalon_rs232_slave_read),       //                   .read
		.write      (mm_interconnect_0_serial_port_avalon_rs232_slave_write),      //                   .write
		.writedata  (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),  //                   .writedata
		.readdata   (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),   //                   .readdata
		.irq        (irq_mapper_receiver5_irq),                                    //          interrupt.irq
		.UART_RXD   (serial_port_external_interface_RXD),                          // external_interface.export
		.UART_TXD   (serial_port_external_interface_TXD)                           //                   .export
	);

	nios_system_sram sram (
		.clk           (sys_clk_out_clk),                                        //                clk.clk
		.reset         (rst_controller_reset_out_reset),                         //              reset.reset
		.SRAM_DQ       (sram_external_interface_DQ),                             // external_interface.export
		.SRAM_ADDR     (sram_external_interface_ADDR),                           //                   .export
		.SRAM_LB_N     (sram_external_interface_LB_N),                           //                   .export
		.SRAM_UB_N     (sram_external_interface_UB_N),                           //                   .export
		.SRAM_CE_N     (sram_external_interface_CE_N),                           //                   .export
		.SRAM_OE_N     (sram_external_interface_OE_N),                           //                   .export
		.SRAM_WE_N     (sram_external_interface_WE_N),                           //                   .export
		.address       (mm_interconnect_0_sram_avalon_sram_slave_address),       //  avalon_sram_slave.address
		.byteenable    (mm_interconnect_0_sram_avalon_sram_slave_byteenable),    //                   .byteenable
		.read          (mm_interconnect_0_sram_avalon_sram_slave_read),          //                   .read
		.write         (mm_interconnect_0_sram_avalon_sram_slave_write),         //                   .write
		.writedata     (mm_interconnect_0_sram_avalon_sram_slave_writedata),     //                   .writedata
		.readdata      (mm_interconnect_0_sram_avalon_sram_slave_readdata),      //                   .readdata
		.readdatavalid (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid)  //                   .readdatavalid
	);

	nios_system_switches switches (
		.clk        (sys_clk_out_clk),                                                  //                        clk.clk
		.reset      (rst_controller_reset_out_reset),                                   //                      reset.reset
		.address    (mm_interconnect_0_switches_avalon_parallel_port_slave_address),    // avalon_parallel_port_slave.address
		.byteenable (mm_interconnect_0_switches_avalon_parallel_port_slave_byteenable), //                           .byteenable
		.chipselect (mm_interconnect_0_switches_avalon_parallel_port_slave_chipselect), //                           .chipselect
		.read       (mm_interconnect_0_switches_avalon_parallel_port_slave_read),       //                           .read
		.write      (mm_interconnect_0_switches_avalon_parallel_port_slave_write),      //                           .write
		.writedata  (mm_interconnect_0_switches_avalon_parallel_port_slave_writedata),  //                           .writedata
		.readdata   (mm_interconnect_0_switches_avalon_parallel_port_slave_readdata),   //                           .readdata
		.SW         (switches_external_interface_export),                               //         external_interface.export
		.irq        (irq_mapper_receiver1_irq)                                          //                  interrupt.irq
	);

	nios_system_sys_sdram_pll sys_sdram_pll (
		.ref_clk_clk        (clk_50_in_clk),                      //      ref_clk.clk
		.ref_reset_reset    (rst_controller_003_reset_out_reset), //    ref_reset.reset
		.sys_clk_clk        (sys_clk_out_clk),                    //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_out_clk),                  //    sdram_clk.clk
		.reset_source_reset (sys_sdram_pll_reset_source_reset)    // reset_source.reset
	);

	nios_system_sysid sysid (
		.clock    (sys_clk_out_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	nios_system_timer timer (
		.clk        (sys_clk_out_clk),                       //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver7_irq)               //   irq.irq
	);

	nios_system_video_chroma_resampler video_chroma_resampler (
		.clk                      (sys_clk_out_clk),                                           //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                            //                reset.reset
		.stream_in_startofpacket  (video_decoder_avalon_decoder_source_startofpacket),         //   avalon_chroma_sink.startofpacket
		.stream_in_endofpacket    (video_decoder_avalon_decoder_source_endofpacket),           //                     .endofpacket
		.stream_in_valid          (video_decoder_avalon_decoder_source_valid),                 //                     .valid
		.stream_in_ready          (video_decoder_avalon_decoder_source_ready),                 //                     .ready
		.stream_in_data           (video_decoder_avalon_decoder_source_data),                  //                     .data
		.stream_out_ready         (video_chroma_resampler_avalon_chroma_source_ready),         // avalon_chroma_source.ready
		.stream_out_startofpacket (video_chroma_resampler_avalon_chroma_source_startofpacket), //                     .startofpacket
		.stream_out_endofpacket   (video_chroma_resampler_avalon_chroma_source_endofpacket),   //                     .endofpacket
		.stream_out_valid         (video_chroma_resampler_avalon_chroma_source_valid),         //                     .valid
		.stream_out_data          (video_chroma_resampler_avalon_chroma_source_data)           //                     .data
	);

	nios_system_video_clipper_normal video_clipper_normal (
		.clk                      (sys_clk_out_clk),                                          //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                           //                 reset.reset
		.stream_in_data           (video_rgb_resampler_avalon_rgb_source_data),               //   avalon_clipper_sink.data
		.stream_in_startofpacket  (video_rgb_resampler_avalon_rgb_source_startofpacket),      //                      .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_avalon_rgb_source_endofpacket),        //                      .endofpacket
		.stream_in_valid          (video_rgb_resampler_avalon_rgb_source_valid),              //                      .valid
		.stream_in_ready          (video_rgb_resampler_avalon_rgb_source_ready),              //                      .ready
		.stream_out_ready         (video_clipper_normal_avalon_clipper_source_ready),         // avalon_clipper_source.ready
		.stream_out_data          (video_clipper_normal_avalon_clipper_source_data),          //                      .data
		.stream_out_startofpacket (video_clipper_normal_avalon_clipper_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_clipper_normal_avalon_clipper_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_clipper_normal_avalon_clipper_source_valid)          //                      .valid
	);

	nios_system_video_csc video_csc (
		.clk                      (sys_clk_out_clk),                                           //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                            //             reset.reset
		.stream_in_startofpacket  (video_chroma_resampler_avalon_chroma_source_startofpacket), //   avalon_csc_sink.startofpacket
		.stream_in_endofpacket    (video_chroma_resampler_avalon_chroma_source_endofpacket),   //                  .endofpacket
		.stream_in_valid          (video_chroma_resampler_avalon_chroma_source_valid),         //                  .valid
		.stream_in_ready          (video_chroma_resampler_avalon_chroma_source_ready),         //                  .ready
		.stream_in_data           (video_chroma_resampler_avalon_chroma_source_data),          //                  .data
		.stream_out_ready         (video_csc_avalon_csc_source_ready),                         // avalon_csc_source.ready
		.stream_out_startofpacket (video_csc_avalon_csc_source_startofpacket),                 //                  .startofpacket
		.stream_out_endofpacket   (video_csc_avalon_csc_source_endofpacket),                   //                  .endofpacket
		.stream_out_valid         (video_csc_avalon_csc_source_valid),                         //                  .valid
		.stream_out_data          (video_csc_avalon_csc_source_data)                           //                  .data
	);

	nios_system_video_decoder video_decoder (
		.clk                      (sys_clk_out_clk),                                   //                   clk.clk
		.reset                    (rst_controller_reset_out_reset),                    //                 reset.reset
		.stream_out_ready         (video_decoder_avalon_decoder_source_ready),         // avalon_decoder_source.ready
		.stream_out_startofpacket (video_decoder_avalon_decoder_source_startofpacket), //                      .startofpacket
		.stream_out_endofpacket   (video_decoder_avalon_decoder_source_endofpacket),   //                      .endofpacket
		.stream_out_valid         (video_decoder_avalon_decoder_source_valid),         //                      .valid
		.stream_out_data          (video_decoder_avalon_decoder_source_data),          //                      .data
		.TD_CLK27                 (video_decoder_external_interface_TD_CLK27),         //    external_interface.export
		.TD_DATA                  (video_decoder_external_interface_TD_DATA),          //                      .export
		.TD_HS                    (video_decoder_external_interface_TD_HS),            //                      .export
		.TD_VS                    (video_decoder_external_interface_TD_VS),            //                      .export
		.clk27_reset              (video_decoder_external_interface_clk27_reset),      //                      .export
		.TD_RESET                 (video_decoder_external_interface_TD_RESET),         //                      .export
		.overflow_flag            (video_decoder_external_interface_overflow_flag)     //                      .export
	);

	nios_system_video_dma_controller_normal video_dma_controller_normal (
		.clk                  (sys_clk_out_clk),                                                                   //                      clk.clk
		.reset                (rst_controller_reset_out_reset),                                                    //                    reset.reset
		.stream_data          (video_scaler_normal_avalon_scaler_source_data),                                     //          avalon_dma_sink.data
		.stream_startofpacket (video_scaler_normal_avalon_scaler_source_startofpacket),                            //                         .startofpacket
		.stream_endofpacket   (video_scaler_normal_avalon_scaler_source_endofpacket),                              //                         .endofpacket
		.stream_valid         (video_scaler_normal_avalon_scaler_source_valid),                                    //                         .valid
		.stream_ready         (video_scaler_normal_avalon_scaler_source_ready),                                    //                         .ready
		.slave_address        (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_address),    // avalon_dma_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_byteenable), //                         .byteenable
		.slave_read           (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_read),       //                         .read
		.slave_write          (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_write),      //                         .write
		.slave_writedata      (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_writedata),  //                         .writedata
		.slave_readdata       (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_readdata),   //                         .readdata
		.master_address       (video_dma_controller_normal_avalon_dma_master_address),                             //        avalon_dma_master.address
		.master_waitrequest   (video_dma_controller_normal_avalon_dma_master_waitrequest),                         //                         .waitrequest
		.master_write         (video_dma_controller_normal_avalon_dma_master_write),                               //                         .write
		.master_writedata     (video_dma_controller_normal_avalon_dma_master_writedata)                            //                         .writedata
	);

	nios_system_video_pll video_pll (
		.ref_clk_clk        (clk_50_2_in_clk),                    //      ref_clk.clk
		.ref_reset_reset    (rst_controller_004_reset_out_reset), //    ref_reset.reset
		.lcd_clk_clk        (mtl_clk_out_clk),                    //      lcd_clk.clk
		.reset_source_reset (video_pll_reset_source_reset)        // reset_source.reset
	);

	nios_system_video_rgb_resampler video_rgb_resampler (
		.clk                      (sys_clk_out_clk),                                     //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                      //             reset.reset
		.stream_in_startofpacket  (video_csc_avalon_csc_source_startofpacket),           //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_csc_avalon_csc_source_endofpacket),             //                  .endofpacket
		.stream_in_valid          (video_csc_avalon_csc_source_valid),                   //                  .valid
		.stream_in_ready          (video_csc_avalon_csc_source_ready),                   //                  .ready
		.stream_in_data           (video_csc_avalon_csc_source_data),                    //                  .data
		.stream_out_ready         (video_rgb_resampler_avalon_rgb_source_ready),         // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_avalon_rgb_source_startofpacket), //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_avalon_rgb_source_endofpacket),   //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_avalon_rgb_source_valid),         //                  .valid
		.stream_out_data          (video_rgb_resampler_avalon_rgb_source_data)           //                  .data
	);

	nios_system_video_scaler_normal video_scaler_normal (
		.clk                      (sys_clk_out_clk),                                          //                  clk.clk
		.reset                    (rst_controller_reset_out_reset),                           //                reset.reset
		.stream_in_startofpacket  (video_clipper_normal_avalon_clipper_source_startofpacket), //   avalon_scaler_sink.startofpacket
		.stream_in_endofpacket    (video_clipper_normal_avalon_clipper_source_endofpacket),   //                     .endofpacket
		.stream_in_valid          (video_clipper_normal_avalon_clipper_source_valid),         //                     .valid
		.stream_in_ready          (video_clipper_normal_avalon_clipper_source_ready),         //                     .ready
		.stream_in_data           (video_clipper_normal_avalon_clipper_source_data),          //                     .data
		.stream_out_ready         (video_scaler_normal_avalon_scaler_source_ready),           // avalon_scaler_source.ready
		.stream_out_startofpacket (video_scaler_normal_avalon_scaler_source_startofpacket),   //                     .startofpacket
		.stream_out_endofpacket   (video_scaler_normal_avalon_scaler_source_endofpacket),     //                     .endofpacket
		.stream_out_valid         (video_scaler_normal_avalon_scaler_source_valid),           //                     .valid
		.stream_out_data          (video_scaler_normal_avalon_scaler_source_data)             //                     .data
	);

	nios_system_mm_interconnect_0 mm_interconnect_0 (
		.sys_sdram_pll_sys_clk_clk                                       (sys_clk_out_clk),                                                                   //                                   sys_sdram_pll_sys_clk.clk
		.video_dma_controller_normal_reset_reset_bridge_in_reset_reset   (rst_controller_reset_out_reset),                                                    // video_dma_controller_normal_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                         (cpu_data_master_address),                                                           //                                         cpu_data_master.address
		.cpu_data_master_waitrequest                                     (cpu_data_master_waitrequest),                                                       //                                                        .waitrequest
		.cpu_data_master_byteenable                                      (cpu_data_master_byteenable),                                                        //                                                        .byteenable
		.cpu_data_master_read                                            (cpu_data_master_read),                                                              //                                                        .read
		.cpu_data_master_readdata                                        (cpu_data_master_readdata),                                                          //                                                        .readdata
		.cpu_data_master_readdatavalid                                   (cpu_data_master_readdatavalid),                                                     //                                                        .readdatavalid
		.cpu_data_master_write                                           (cpu_data_master_write),                                                             //                                                        .write
		.cpu_data_master_writedata                                       (cpu_data_master_writedata),                                                         //                                                        .writedata
		.cpu_data_master_debugaccess                                     (cpu_data_master_debugaccess),                                                       //                                                        .debugaccess
		.cpu_instruction_master_address                                  (cpu_instruction_master_address),                                                    //                                  cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                              (cpu_instruction_master_waitrequest),                                                //                                                        .waitrequest
		.cpu_instruction_master_read                                     (cpu_instruction_master_read),                                                       //                                                        .read
		.cpu_instruction_master_readdata                                 (cpu_instruction_master_readdata),                                                   //                                                        .readdata
		.cpu_instruction_master_readdatavalid                            (cpu_instruction_master_readdatavalid),                                              //                                                        .readdatavalid
		.pixel_buffer_dma_green_avalon_pixel_dma_master_address          (pixel_buffer_dma_green_avalon_pixel_dma_master_address),                            //          pixel_buffer_dma_green_avalon_pixel_dma_master.address
		.pixel_buffer_dma_green_avalon_pixel_dma_master_waitrequest      (pixel_buffer_dma_green_avalon_pixel_dma_master_waitrequest),                        //                                                        .waitrequest
		.pixel_buffer_dma_green_avalon_pixel_dma_master_read             (pixel_buffer_dma_green_avalon_pixel_dma_master_read),                               //                                                        .read
		.pixel_buffer_dma_green_avalon_pixel_dma_master_readdata         (pixel_buffer_dma_green_avalon_pixel_dma_master_readdata),                           //                                                        .readdata
		.pixel_buffer_dma_green_avalon_pixel_dma_master_readdatavalid    (pixel_buffer_dma_green_avalon_pixel_dma_master_readdatavalid),                      //                                                        .readdatavalid
		.pixel_buffer_dma_green_avalon_pixel_dma_master_lock             (pixel_buffer_dma_green_avalon_pixel_dma_master_lock),                               //                                                        .lock
		.video_dma_controller_normal_avalon_dma_master_address           (video_dma_controller_normal_avalon_dma_master_address),                             //           video_dma_controller_normal_avalon_dma_master.address
		.video_dma_controller_normal_avalon_dma_master_waitrequest       (video_dma_controller_normal_avalon_dma_master_waitrequest),                         //                                                        .waitrequest
		.video_dma_controller_normal_avalon_dma_master_write             (video_dma_controller_normal_avalon_dma_master_write),                               //                                                        .write
		.video_dma_controller_normal_avalon_dma_master_writedata         (video_dma_controller_normal_avalon_dma_master_writedata),                           //                                                        .writedata
		.audio_avalon_audio_slave_address                                (mm_interconnect_0_audio_avalon_audio_slave_address),                                //                                audio_avalon_audio_slave.address
		.audio_avalon_audio_slave_write                                  (mm_interconnect_0_audio_avalon_audio_slave_write),                                  //                                                        .write
		.audio_avalon_audio_slave_read                                   (mm_interconnect_0_audio_avalon_audio_slave_read),                                   //                                                        .read
		.audio_avalon_audio_slave_readdata                               (mm_interconnect_0_audio_avalon_audio_slave_readdata),                               //                                                        .readdata
		.audio_avalon_audio_slave_writedata                              (mm_interconnect_0_audio_avalon_audio_slave_writedata),                              //                                                        .writedata
		.audio_avalon_audio_slave_chipselect                             (mm_interconnect_0_audio_avalon_audio_slave_chipselect),                             //                                                        .chipselect
		.audio_and_video_config_avalon_av_config_slave_address           (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_address),           //           audio_and_video_config_avalon_av_config_slave.address
		.audio_and_video_config_avalon_av_config_slave_write             (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_write),             //                                                        .write
		.audio_and_video_config_avalon_av_config_slave_read              (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_read),              //                                                        .read
		.audio_and_video_config_avalon_av_config_slave_readdata          (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_readdata),          //                                                        .readdata
		.audio_and_video_config_avalon_av_config_slave_writedata         (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_writedata),         //                                                        .writedata
		.audio_and_video_config_avalon_av_config_slave_byteenable        (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_byteenable),        //                                                        .byteenable
		.audio_and_video_config_avalon_av_config_slave_waitrequest       (mm_interconnect_0_audio_and_video_config_avalon_av_config_slave_waitrequest),       //                                                        .waitrequest
		.char_lcd_avalon_lcd_slave_address                               (mm_interconnect_0_char_lcd_avalon_lcd_slave_address),                               //                               char_lcd_avalon_lcd_slave.address
		.char_lcd_avalon_lcd_slave_write                                 (mm_interconnect_0_char_lcd_avalon_lcd_slave_write),                                 //                                                        .write
		.char_lcd_avalon_lcd_slave_read                                  (mm_interconnect_0_char_lcd_avalon_lcd_slave_read),                                  //                                                        .read
		.char_lcd_avalon_lcd_slave_readdata                              (mm_interconnect_0_char_lcd_avalon_lcd_slave_readdata),                              //                                                        .readdata
		.char_lcd_avalon_lcd_slave_writedata                             (mm_interconnect_0_char_lcd_avalon_lcd_slave_writedata),                             //                                                        .writedata
		.char_lcd_avalon_lcd_slave_waitrequest                           (mm_interconnect_0_char_lcd_avalon_lcd_slave_waitrequest),                           //                                                        .waitrequest
		.char_lcd_avalon_lcd_slave_chipselect                            (mm_interconnect_0_char_lcd_avalon_lcd_slave_chipselect),                            //                                                        .chipselect
		.cpu_debug_mem_slave_address                                     (mm_interconnect_0_cpu_debug_mem_slave_address),                                     //                                     cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                                       (mm_interconnect_0_cpu_debug_mem_slave_write),                                       //                                                        .write
		.cpu_debug_mem_slave_read                                        (mm_interconnect_0_cpu_debug_mem_slave_read),                                        //                                                        .read
		.cpu_debug_mem_slave_readdata                                    (mm_interconnect_0_cpu_debug_mem_slave_readdata),                                    //                                                        .readdata
		.cpu_debug_mem_slave_writedata                                   (mm_interconnect_0_cpu_debug_mem_slave_writedata),                                   //                                                        .writedata
		.cpu_debug_mem_slave_byteenable                                  (mm_interconnect_0_cpu_debug_mem_slave_byteenable),                                  //                                                        .byteenable
		.cpu_debug_mem_slave_waitrequest                                 (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),                                 //                                                        .waitrequest
		.cpu_debug_mem_slave_debugaccess                                 (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),                                 //                                                        .debugaccess
		.flash_controller_uas_address                                    (mm_interconnect_0_flash_controller_uas_address),                                    //                                    flash_controller_uas.address
		.flash_controller_uas_write                                      (mm_interconnect_0_flash_controller_uas_write),                                      //                                                        .write
		.flash_controller_uas_read                                       (mm_interconnect_0_flash_controller_uas_read),                                       //                                                        .read
		.flash_controller_uas_readdata                                   (mm_interconnect_0_flash_controller_uas_readdata),                                   //                                                        .readdata
		.flash_controller_uas_writedata                                  (mm_interconnect_0_flash_controller_uas_writedata),                                  //                                                        .writedata
		.flash_controller_uas_burstcount                                 (mm_interconnect_0_flash_controller_uas_burstcount),                                 //                                                        .burstcount
		.flash_controller_uas_byteenable                                 (mm_interconnect_0_flash_controller_uas_byteenable),                                 //                                                        .byteenable
		.flash_controller_uas_readdatavalid                              (mm_interconnect_0_flash_controller_uas_readdatavalid),                              //                                                        .readdatavalid
		.flash_controller_uas_waitrequest                                (mm_interconnect_0_flash_controller_uas_waitrequest),                                //                                                        .waitrequest
		.flash_controller_uas_lock                                       (mm_interconnect_0_flash_controller_uas_lock),                                       //                                                        .lock
		.flash_controller_uas_debugaccess                                (mm_interconnect_0_flash_controller_uas_debugaccess),                                //                                                        .debugaccess
		.Green_LED_avalon_parallel_port_slave_address                    (mm_interconnect_0_green_led_avalon_parallel_port_slave_address),                    //                    Green_LED_avalon_parallel_port_slave.address
		.Green_LED_avalon_parallel_port_slave_write                      (mm_interconnect_0_green_led_avalon_parallel_port_slave_write),                      //                                                        .write
		.Green_LED_avalon_parallel_port_slave_read                       (mm_interconnect_0_green_led_avalon_parallel_port_slave_read),                       //                                                        .read
		.Green_LED_avalon_parallel_port_slave_readdata                   (mm_interconnect_0_green_led_avalon_parallel_port_slave_readdata),                   //                                                        .readdata
		.Green_LED_avalon_parallel_port_slave_writedata                  (mm_interconnect_0_green_led_avalon_parallel_port_slave_writedata),                  //                                                        .writedata
		.Green_LED_avalon_parallel_port_slave_byteenable                 (mm_interconnect_0_green_led_avalon_parallel_port_slave_byteenable),                 //                                                        .byteenable
		.Green_LED_avalon_parallel_port_slave_chipselect                 (mm_interconnect_0_green_led_avalon_parallel_port_slave_chipselect),                 //                                                        .chipselect
		.HEX3_HEX0_avalon_parallel_port_slave_address                    (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_address),                    //                    HEX3_HEX0_avalon_parallel_port_slave.address
		.HEX3_HEX0_avalon_parallel_port_slave_write                      (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_write),                      //                                                        .write
		.HEX3_HEX0_avalon_parallel_port_slave_read                       (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_read),                       //                                                        .read
		.HEX3_HEX0_avalon_parallel_port_slave_readdata                   (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_readdata),                   //                                                        .readdata
		.HEX3_HEX0_avalon_parallel_port_slave_writedata                  (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_writedata),                  //                                                        .writedata
		.HEX3_HEX0_avalon_parallel_port_slave_byteenable                 (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_byteenable),                 //                                                        .byteenable
		.HEX3_HEX0_avalon_parallel_port_slave_chipselect                 (mm_interconnect_0_hex3_hex0_avalon_parallel_port_slave_chipselect),                 //                                                        .chipselect
		.HEX7_HEX4_avalon_parallel_port_slave_address                    (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_address),                    //                    HEX7_HEX4_avalon_parallel_port_slave.address
		.HEX7_HEX4_avalon_parallel_port_slave_write                      (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_write),                      //                                                        .write
		.HEX7_HEX4_avalon_parallel_port_slave_read                       (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_read),                       //                                                        .read
		.HEX7_HEX4_avalon_parallel_port_slave_readdata                   (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_readdata),                   //                                                        .readdata
		.HEX7_HEX4_avalon_parallel_port_slave_writedata                  (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_writedata),                  //                                                        .writedata
		.HEX7_HEX4_avalon_parallel_port_slave_byteenable                 (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_byteenable),                 //                                                        .byteenable
		.HEX7_HEX4_avalon_parallel_port_slave_chipselect                 (mm_interconnect_0_hex7_hex4_avalon_parallel_port_slave_chipselect),                 //                                                        .chipselect
		.jtag_uart_avalon_jtag_slave_address                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),                             //                             jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),                               //                                                        .write
		.jtag_uart_avalon_jtag_slave_read                                (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),                                //                                                        .read
		.jtag_uart_avalon_jtag_slave_readdata                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),                            //                                                        .readdata
		.jtag_uart_avalon_jtag_slave_writedata                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),                           //                                                        .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),                         //                                                        .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),                          //                                                        .chipselect
		.mtl_char_buffer_avalon_char_buffer_slave_address                (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_address),                //                mtl_char_buffer_avalon_char_buffer_slave.address
		.mtl_char_buffer_avalon_char_buffer_slave_write                  (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_write),                  //                                                        .write
		.mtl_char_buffer_avalon_char_buffer_slave_read                   (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_read),                   //                                                        .read
		.mtl_char_buffer_avalon_char_buffer_slave_readdata               (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_readdata),               //                                                        .readdata
		.mtl_char_buffer_avalon_char_buffer_slave_writedata              (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_writedata),              //                                                        .writedata
		.mtl_char_buffer_avalon_char_buffer_slave_byteenable             (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_byteenable),             //                                                        .byteenable
		.mtl_char_buffer_avalon_char_buffer_slave_waitrequest            (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_waitrequest),            //                                                        .waitrequest
		.mtl_char_buffer_avalon_char_buffer_slave_chipselect             (mm_interconnect_0_mtl_char_buffer_avalon_char_buffer_slave_chipselect),             //                                                        .chipselect
		.mtl_char_buffer_avalon_char_control_slave_address               (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_address),               //               mtl_char_buffer_avalon_char_control_slave.address
		.mtl_char_buffer_avalon_char_control_slave_write                 (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_write),                 //                                                        .write
		.mtl_char_buffer_avalon_char_control_slave_read                  (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_read),                  //                                                        .read
		.mtl_char_buffer_avalon_char_control_slave_readdata              (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_readdata),              //                                                        .readdata
		.mtl_char_buffer_avalon_char_control_slave_writedata             (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_writedata),             //                                                        .writedata
		.mtl_char_buffer_avalon_char_control_slave_byteenable            (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_byteenable),            //                                                        .byteenable
		.mtl_char_buffer_avalon_char_control_slave_chipselect            (mm_interconnect_0_mtl_char_buffer_avalon_char_control_slave_chipselect),            //                                                        .chipselect
		.onchip_memory_s1_address                                        (mm_interconnect_0_onchip_memory_s1_address),                                        //                                        onchip_memory_s1.address
		.onchip_memory_s1_write                                          (mm_interconnect_0_onchip_memory_s1_write),                                          //                                                        .write
		.onchip_memory_s1_readdata                                       (mm_interconnect_0_onchip_memory_s1_readdata),                                       //                                                        .readdata
		.onchip_memory_s1_writedata                                      (mm_interconnect_0_onchip_memory_s1_writedata),                                      //                                                        .writedata
		.onchip_memory_s1_byteenable                                     (mm_interconnect_0_onchip_memory_s1_byteenable),                                     //                                                        .byteenable
		.onchip_memory_s1_chipselect                                     (mm_interconnect_0_onchip_memory_s1_chipselect),                                     //                                                        .chipselect
		.onchip_memory_s1_clken                                          (mm_interconnect_0_onchip_memory_s1_clken),                                          //                                                        .clken
		.performance_counter_control_slave_address                       (mm_interconnect_0_performance_counter_control_slave_address),                       //                       performance_counter_control_slave.address
		.performance_counter_control_slave_write                         (mm_interconnect_0_performance_counter_control_slave_write),                         //                                                        .write
		.performance_counter_control_slave_readdata                      (mm_interconnect_0_performance_counter_control_slave_readdata),                      //                                                        .readdata
		.performance_counter_control_slave_writedata                     (mm_interconnect_0_performance_counter_control_slave_writedata),                     //                                                        .writedata
		.performance_counter_control_slave_begintransfer                 (mm_interconnect_0_performance_counter_control_slave_begintransfer),                 //                                                        .begintransfer
		.pixel_buffer_dma_green_avalon_control_slave_address             (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_address),             //             pixel_buffer_dma_green_avalon_control_slave.address
		.pixel_buffer_dma_green_avalon_control_slave_write               (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_write),               //                                                        .write
		.pixel_buffer_dma_green_avalon_control_slave_read                (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_read),                //                                                        .read
		.pixel_buffer_dma_green_avalon_control_slave_readdata            (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_readdata),            //                                                        .readdata
		.pixel_buffer_dma_green_avalon_control_slave_writedata           (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_writedata),           //                                                        .writedata
		.pixel_buffer_dma_green_avalon_control_slave_byteenable          (mm_interconnect_0_pixel_buffer_dma_green_avalon_control_slave_byteenable),          //                                                        .byteenable
		.ps2_key_avalon_ps2_slave_address                                (mm_interconnect_0_ps2_key_avalon_ps2_slave_address),                                //                                ps2_key_avalon_ps2_slave.address
		.ps2_key_avalon_ps2_slave_write                                  (mm_interconnect_0_ps2_key_avalon_ps2_slave_write),                                  //                                                        .write
		.ps2_key_avalon_ps2_slave_read                                   (mm_interconnect_0_ps2_key_avalon_ps2_slave_read),                                   //                                                        .read
		.ps2_key_avalon_ps2_slave_readdata                               (mm_interconnect_0_ps2_key_avalon_ps2_slave_readdata),                               //                                                        .readdata
		.ps2_key_avalon_ps2_slave_writedata                              (mm_interconnect_0_ps2_key_avalon_ps2_slave_writedata),                              //                                                        .writedata
		.ps2_key_avalon_ps2_slave_byteenable                             (mm_interconnect_0_ps2_key_avalon_ps2_slave_byteenable),                             //                                                        .byteenable
		.ps2_key_avalon_ps2_slave_waitrequest                            (mm_interconnect_0_ps2_key_avalon_ps2_slave_waitrequest),                            //                                                        .waitrequest
		.ps2_key_avalon_ps2_slave_chipselect                             (mm_interconnect_0_ps2_key_avalon_ps2_slave_chipselect),                             //                                                        .chipselect
		.ps2_mouse_avalon_ps2_slave_address                              (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_address),                              //                              ps2_mouse_avalon_ps2_slave.address
		.ps2_mouse_avalon_ps2_slave_write                                (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_write),                                //                                                        .write
		.ps2_mouse_avalon_ps2_slave_read                                 (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_read),                                 //                                                        .read
		.ps2_mouse_avalon_ps2_slave_readdata                             (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_readdata),                             //                                                        .readdata
		.ps2_mouse_avalon_ps2_slave_writedata                            (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_writedata),                            //                                                        .writedata
		.ps2_mouse_avalon_ps2_slave_byteenable                           (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_byteenable),                           //                                                        .byteenable
		.ps2_mouse_avalon_ps2_slave_waitrequest                          (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_waitrequest),                          //                                                        .waitrequest
		.ps2_mouse_avalon_ps2_slave_chipselect                           (mm_interconnect_0_ps2_mouse_avalon_ps2_slave_chipselect),                           //                                                        .chipselect
		.pushbuttons_avalon_parallel_port_slave_address                  (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_address),                  //                  pushbuttons_avalon_parallel_port_slave.address
		.pushbuttons_avalon_parallel_port_slave_write                    (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_write),                    //                                                        .write
		.pushbuttons_avalon_parallel_port_slave_read                     (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_read),                     //                                                        .read
		.pushbuttons_avalon_parallel_port_slave_readdata                 (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_readdata),                 //                                                        .readdata
		.pushbuttons_avalon_parallel_port_slave_writedata                (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_writedata),                //                                                        .writedata
		.pushbuttons_avalon_parallel_port_slave_byteenable               (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_byteenable),               //                                                        .byteenable
		.pushbuttons_avalon_parallel_port_slave_chipselect               (mm_interconnect_0_pushbuttons_avalon_parallel_port_slave_chipselect),               //                                                        .chipselect
		.red_LEDs_avalon_parallel_port_slave_address                     (mm_interconnect_0_red_leds_avalon_parallel_port_slave_address),                     //                     red_LEDs_avalon_parallel_port_slave.address
		.red_LEDs_avalon_parallel_port_slave_write                       (mm_interconnect_0_red_leds_avalon_parallel_port_slave_write),                       //                                                        .write
		.red_LEDs_avalon_parallel_port_slave_read                        (mm_interconnect_0_red_leds_avalon_parallel_port_slave_read),                        //                                                        .read
		.red_LEDs_avalon_parallel_port_slave_readdata                    (mm_interconnect_0_red_leds_avalon_parallel_port_slave_readdata),                    //                                                        .readdata
		.red_LEDs_avalon_parallel_port_slave_writedata                   (mm_interconnect_0_red_leds_avalon_parallel_port_slave_writedata),                   //                                                        .writedata
		.red_LEDs_avalon_parallel_port_slave_byteenable                  (mm_interconnect_0_red_leds_avalon_parallel_port_slave_byteenable),                  //                                                        .byteenable
		.red_LEDs_avalon_parallel_port_slave_chipselect                  (mm_interconnect_0_red_leds_avalon_parallel_port_slave_chipselect),                  //                                                        .chipselect
		.sd_card_avalon_sdcard_slave_address                             (mm_interconnect_0_sd_card_avalon_sdcard_slave_address),                             //                             sd_card_avalon_sdcard_slave.address
		.sd_card_avalon_sdcard_slave_write                               (mm_interconnect_0_sd_card_avalon_sdcard_slave_write),                               //                                                        .write
		.sd_card_avalon_sdcard_slave_read                                (mm_interconnect_0_sd_card_avalon_sdcard_slave_read),                                //                                                        .read
		.sd_card_avalon_sdcard_slave_readdata                            (mm_interconnect_0_sd_card_avalon_sdcard_slave_readdata),                            //                                                        .readdata
		.sd_card_avalon_sdcard_slave_writedata                           (mm_interconnect_0_sd_card_avalon_sdcard_slave_writedata),                           //                                                        .writedata
		.sd_card_avalon_sdcard_slave_byteenable                          (mm_interconnect_0_sd_card_avalon_sdcard_slave_byteenable),                          //                                                        .byteenable
		.sd_card_avalon_sdcard_slave_waitrequest                         (mm_interconnect_0_sd_card_avalon_sdcard_slave_waitrequest),                         //                                                        .waitrequest
		.sd_card_avalon_sdcard_slave_chipselect                          (mm_interconnect_0_sd_card_avalon_sdcard_slave_chipselect),                          //                                                        .chipselect
		.sdram_s1_address                                                (mm_interconnect_0_sdram_s1_address),                                                //                                                sdram_s1.address
		.sdram_s1_write                                                  (mm_interconnect_0_sdram_s1_write),                                                  //                                                        .write
		.sdram_s1_read                                                   (mm_interconnect_0_sdram_s1_read),                                                   //                                                        .read
		.sdram_s1_readdata                                               (mm_interconnect_0_sdram_s1_readdata),                                               //                                                        .readdata
		.sdram_s1_writedata                                              (mm_interconnect_0_sdram_s1_writedata),                                              //                                                        .writedata
		.sdram_s1_byteenable                                             (mm_interconnect_0_sdram_s1_byteenable),                                             //                                                        .byteenable
		.sdram_s1_readdatavalid                                          (mm_interconnect_0_sdram_s1_readdatavalid),                                          //                                                        .readdatavalid
		.sdram_s1_waitrequest                                            (mm_interconnect_0_sdram_s1_waitrequest),                                            //                                                        .waitrequest
		.sdram_s1_chipselect                                             (mm_interconnect_0_sdram_s1_chipselect),                                             //                                                        .chipselect
		.serial_port_avalon_rs232_slave_address                          (mm_interconnect_0_serial_port_avalon_rs232_slave_address),                          //                          serial_port_avalon_rs232_slave.address
		.serial_port_avalon_rs232_slave_write                            (mm_interconnect_0_serial_port_avalon_rs232_slave_write),                            //                                                        .write
		.serial_port_avalon_rs232_slave_read                             (mm_interconnect_0_serial_port_avalon_rs232_slave_read),                             //                                                        .read
		.serial_port_avalon_rs232_slave_readdata                         (mm_interconnect_0_serial_port_avalon_rs232_slave_readdata),                         //                                                        .readdata
		.serial_port_avalon_rs232_slave_writedata                        (mm_interconnect_0_serial_port_avalon_rs232_slave_writedata),                        //                                                        .writedata
		.serial_port_avalon_rs232_slave_byteenable                       (mm_interconnect_0_serial_port_avalon_rs232_slave_byteenable),                       //                                                        .byteenable
		.serial_port_avalon_rs232_slave_chipselect                       (mm_interconnect_0_serial_port_avalon_rs232_slave_chipselect),                       //                                                        .chipselect
		.sram_avalon_sram_slave_address                                  (mm_interconnect_0_sram_avalon_sram_slave_address),                                  //                                  sram_avalon_sram_slave.address
		.sram_avalon_sram_slave_write                                    (mm_interconnect_0_sram_avalon_sram_slave_write),                                    //                                                        .write
		.sram_avalon_sram_slave_read                                     (mm_interconnect_0_sram_avalon_sram_slave_read),                                     //                                                        .read
		.sram_avalon_sram_slave_readdata                                 (mm_interconnect_0_sram_avalon_sram_slave_readdata),                                 //                                                        .readdata
		.sram_avalon_sram_slave_writedata                                (mm_interconnect_0_sram_avalon_sram_slave_writedata),                                //                                                        .writedata
		.sram_avalon_sram_slave_byteenable                               (mm_interconnect_0_sram_avalon_sram_slave_byteenable),                               //                                                        .byteenable
		.sram_avalon_sram_slave_readdatavalid                            (mm_interconnect_0_sram_avalon_sram_slave_readdatavalid),                            //                                                        .readdatavalid
		.switches_avalon_parallel_port_slave_address                     (mm_interconnect_0_switches_avalon_parallel_port_slave_address),                     //                     switches_avalon_parallel_port_slave.address
		.switches_avalon_parallel_port_slave_write                       (mm_interconnect_0_switches_avalon_parallel_port_slave_write),                       //                                                        .write
		.switches_avalon_parallel_port_slave_read                        (mm_interconnect_0_switches_avalon_parallel_port_slave_read),                        //                                                        .read
		.switches_avalon_parallel_port_slave_readdata                    (mm_interconnect_0_switches_avalon_parallel_port_slave_readdata),                    //                                                        .readdata
		.switches_avalon_parallel_port_slave_writedata                   (mm_interconnect_0_switches_avalon_parallel_port_slave_writedata),                   //                                                        .writedata
		.switches_avalon_parallel_port_slave_byteenable                  (mm_interconnect_0_switches_avalon_parallel_port_slave_byteenable),                  //                                                        .byteenable
		.switches_avalon_parallel_port_slave_chipselect                  (mm_interconnect_0_switches_avalon_parallel_port_slave_chipselect),                  //                                                        .chipselect
		.sysid_control_slave_address                                     (mm_interconnect_0_sysid_control_slave_address),                                     //                                     sysid_control_slave.address
		.sysid_control_slave_readdata                                    (mm_interconnect_0_sysid_control_slave_readdata),                                    //                                                        .readdata
		.timer_s1_address                                                (mm_interconnect_0_timer_s1_address),                                                //                                                timer_s1.address
		.timer_s1_write                                                  (mm_interconnect_0_timer_s1_write),                                                  //                                                        .write
		.timer_s1_readdata                                               (mm_interconnect_0_timer_s1_readdata),                                               //                                                        .readdata
		.timer_s1_writedata                                              (mm_interconnect_0_timer_s1_writedata),                                              //                                                        .writedata
		.timer_s1_chipselect                                             (mm_interconnect_0_timer_s1_chipselect),                                             //                                                        .chipselect
		.video_dma_controller_normal_avalon_dma_control_slave_address    (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_address),    //    video_dma_controller_normal_avalon_dma_control_slave.address
		.video_dma_controller_normal_avalon_dma_control_slave_write      (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_write),      //                                                        .write
		.video_dma_controller_normal_avalon_dma_control_slave_read       (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_read),       //                                                        .read
		.video_dma_controller_normal_avalon_dma_control_slave_readdata   (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_readdata),   //                                                        .readdata
		.video_dma_controller_normal_avalon_dma_control_slave_writedata  (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_writedata),  //                                                        .writedata
		.video_dma_controller_normal_avalon_dma_control_slave_byteenable (mm_interconnect_0_video_dma_controller_normal_avalon_dma_control_slave_byteenable)  //                                                        .byteenable
	);

	nios_system_irq_mapper irq_mapper (
		.clk           (sys_clk_out_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),       // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),       // receiver7.irq
		.sender_irq    (cpu_irq_irq)                     //    sender.irq
	);

	nios_system_avalon_st_adapter #(
		.inBitsPerSymbol (10),
		.inUsePackets    (1),
		.inDataWidth     (30),
		.inChannelWidth  (2),
		.inErrorWidth    (0),
		.inUseEmptyPort  (0),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (0),
		.outDataWidth    (30),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (sys_clk_out_clk),                                 // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_reset_out_reset),                  // in_rst_0.reset
		.in_0_data           (scaler_green_avalon_scaler_source_data),          //     in_0.data
		.in_0_valid          (scaler_green_avalon_scaler_source_valid),         //         .valid
		.in_0_ready          (scaler_green_avalon_scaler_source_ready),         //         .ready
		.in_0_startofpacket  (scaler_green_avalon_scaler_source_startofpacket), //         .startofpacket
		.in_0_endofpacket    (scaler_green_avalon_scaler_source_endofpacket),   //         .endofpacket
		.in_0_channel        (scaler_green_avalon_scaler_source_channel),       //         .channel
		.out_0_data          (avalon_st_adapter_out_0_data),                    //    out_0.data
		.out_0_valid         (avalon_st_adapter_out_0_valid),                   //         .valid
		.out_0_ready         (avalon_st_adapter_out_0_ready),                   //         .ready
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket),           //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)              //         .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (sys_sdram_pll_reset_source_reset),   // reset_in1.reset
		.clk            (sys_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_bridge_in_reset_n),           // reset_in0.reset
		.clk            (clk_50_3_in_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_debug_reset_request_reset),      // reset_in0.reset
		.reset_in1      (video_pll_reset_source_reset),       // reset_in1.reset
		.clk            (mtl_clk_out_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_bridge_in_reset_n),           // reset_in0.reset
		.clk            (clk_50_in_clk),                      //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_bridge_in_reset_n),           // reset_in0.reset
		.clk            (clk_50_2_in_clk),                    //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
